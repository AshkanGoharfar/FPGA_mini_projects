`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
qbPtSB0hCgD8MlHzYH3+RfAdhQfC6Jls3IexjyuBIVvModTNrehm1/fydUmgQwgzWFu5ePOpAroW
mjAP232h7Q==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
HO57n6yJr04IaE3Mpu434kjt8GjGB0Hi2pvizhtf/BH1RvBygoGQSNk9h+sHAQDQxe09pbpCq77W
ThmIuMfzSZKOi/tOo6dcHmCJVpdgaNH2qjSYNdKy4x8biS38ihYMKcGImLqxrDD4UKPaxV2Ef16L
jtajkQUbyke0nxKsyc4=

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
rLgwFZ3dPgt8Q5fdSWPl0ix9QMgOtsTUT8bQR5EfrmAmMrpF7IHR3gKNzq18SCY3H8+AznDiesny
i32h5U2ZtUHf5qtVyJx56jGgMkeo7ylXXIVnEuNSVEggRRgwFewddWXDf+Ol7iF8jwWfGVUHDcRJ
FEJQpejowcye/lCCE6Q=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
XQUH5+FuZVQ/kTB2wgYB8j8qARHhWqWb0NV6dEttAxL2q3VyoNg14pl6VWP7QW3yGvJctKo7PZDW
bhc2cO+h5vUaOjPgT6u9wEUbMxtMROV+KnEbvv3QOMYyxz792eY2Hsy/3QG33+3yXJkTVh88xNUa
+nzcfXtBe+TFmX/jzy/q1mV47vmki8Mzcst9EAkfk6Ewjn5z98/5DOqUUUTWS3fG5E8AZLWKD76h
nuOh9sc04HFc8TZvxjRy2xbmJa+cQjM7QBvigGdd6k1fwjEvn+OpNywKd3rBXdk0tGZSppIf04Lz
fzDHI/4hV7KBDAeAc68yu4NOHFK5umSC5TXjLg==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
P5jOSAc+0BlAfnLcoWZLfuF/cUc8LfYQspxB1Jha/9RAHr0cCXkFeGwBmzKHPOUllv73ghBuPnZW
Qnky4ctPauhdPSlgBVhEK3oDBriwkG/nhI3BMwI9Z5BNByJ7Mrr0eD6sR0gYWkTg/vbUYeSA6FI4
RBpTxspkssZ7GrD1TGxn348ZZL5Z5onGFZ+Lq7SSRacXPtU83RtCSs1rREXpMeueCWxYxJ0+uzwc
WRtWTUWIkSzfcvgKSobhmWhAyogWNaNZkBfh5STy7d3mj1/UF7XOuycrSW1a5va7agOibrEbbXh9
4pdS6h+61DPvePev9unaTBCvHqGvYt+gewy4Cw==

`protect key_keyowner = "Xilinx", key_keyname = "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
rtGfi6/RX0wsETsRTgqAqouM8WkNinF3NEq+iUVhGe1BgHYmE369Eqa/qMqePosSehXlvcQt9vhe
d1GgGf/hfbIaGGa+YjleJNpbaj7v3jXX9C7y2g8B1ji018c2JRlFIfSpiXArfhl3GiZblSgfqDW1
/iq01P0SR5QNlyIVLhxOnLD4bD3nx4jt6zzbVCHmv0CRMokD8AuI+I2lDpPzHgwFzcPwh7fCqpBX
4xU6Nd2Qs3bJzKE2tHy/Uo0j0mCjaOQlRhvCKVE++p8Kp58TTknYaLUhvj9sEb+aQXsqH8fAjqqK
cBCpAgZjBeK2ap16L8lpjSdKnUC8rmBMaoVdPA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 63104)
`protect data_block
0J4NlSx8TF5s82HxqudqKtK3SE5NP1zOq2ULJQhzOBaqZ4KzFz+w6NZljnValemx5WutVYzUbIdY
WD835PSj+8X86NdZYdDn2a+jDzmd6wZf8sFU6qFqHUF1yaIBy+p+W8ELaQ+1WdLZzNxZTR6Tc85m
Fa5Js5XsfriGm06efgrCNj3tV2pFOKtc8nmuIy/9wxy0RPx7jrAaHaz9ChU+0nCPGvtzCIxMR24y
RD3LUY+o/gw6rkVEafI0XsNTKiP5ADXxihH3MAmStMTZSW5OwMjRIO5jawbSH3Laa6KkW0SHaEph
1y467KxYidPT6Q1tYQ/lpqCDeQ47UTr8GcheEPJJ3h47h0aOgP6Lz/4CuhUOHWpHw/lBnxNX40wD
V8xzv+Od0fSXR6SDGURgg82MlOpUSgYBaqHqiuYBYkVJLspFgDeXQEU5Pj9s1m5iS3p9ViLVs6Xi
5pAZ5XQipaWhmBc23SqoBctc+6xKsu8Y0hqlEZ3hl69r3pOOG+Bo5qG+jgWbxRS9sdJdDiU1sXCG
fqI4pOi/QLm/2kAlLv0x+U+FFXt1Gt2kqSe//1fyf1d/lN5PeKfC7h+z9ibRYbc/DjMP9aYmrpR3
wfFG5R8ap3jlOScins/GDT78np3EF3Hl8eEFiVbad13F7VUEs/AjSrzYv/IOYTARwWguPkfnos2U
A4ySx2ILVTa7VuWYG7T1ILPIwe1tNn+ok24XSeCAuLmqqVmev08fLIt04HD892EdfsPHSSaoXrZr
cWT3KNtySHZddvc5/o175AGdZ6wf0q1TFBO+N9GU/zW7jmNwWSOFIkcNzqvwAng53zKz8mFuAMGq
zaW30frMGeSqg/E67dSVX/0PUJNhjo+eWWnfdZm6nLrFdU0hDsF4hZPBydanxg7gijflGc4UFjUR
eyZbWkVUpQMCRt7xnhR3qwSKilvPmXYOgye+/NZvgdteHlCUl6ies9/owPypfAg2svajjXn9RKYk
kjFbdlRhikxfQo9nQq+oBDYetGBcZ/0jvcheGGO4T7FKgnM1Clnnq1NWeUosegdI8z9630wvL54C
T5ELYant1C5+R2vxsYrbVtGemASYiYjbkbRuw2jkQvVJq2Y4DdVEEc53+5GxtPP8EKpjO38hyIX2
8YWl3g/sDOCYWoRW4H3hc4XXUAlYNUZtF+z2VjUB9bqlR9V2/3ehiHMqAtvfbDKv1USIzw4wdF9o
C/4wfo21PxjJYmoRqL7T5ycDRDafrN3DKWAw2X70HPtejpkJ8SYdyZFvzrA5y/LybuthGqs8uKlu
VNnd/pKBl1slEuGMVgqUJ06KnwmbaPvv5JVR3sLMJnMGoKA8vuwMdXkBKSLhkh2Tw2PkowbkYwVd
cmTL69HxZfOhBRKZXO+rFRr2yGLUzZ0mlMqONUF6KVejJMOhX3tSKy3KjM+T42Tgj8+MUBgGbx8j
1sojPwQXIU1SN8M6atU1rSTTLuJXaN48C3xXZA1bSfR27iI+ygIKgPE8PWQFSKHvL+IaUPELLtJk
pmKBmbSq86/xvYrvUpLvFrGogHVd1pyWAPDxpNjF+Fq75FFV/7wGo0M+eHGHRpLhEwpuSmxIfF1C
FDXu2rBmYHvuu0zaWNH8CGf09pFvEi7nf46zuAheF/sYdpJQJkCkDDmE3CcLFLhjTXcVwCyurhic
I1Y7mmeHF+vU5ZzMm2dk+hxQzZehaShaDmLTVPifgHhXYg4HBB5seeaJRLpsqW3gbFhsJxYVbwfi
F2MwEH9Xd3ehj2YRYi4tgExtceRTF7ArfoYYmW1a5+s8J+WZU4Cxh+AUQA+nC6wG4F5fSdTY4mEo
pvIt7UvAXCDbaytLVi7Cgh+BLvJRWT4bO1hNxO1oLjdjihY4SsGkN8OgVgdur2jLWZtd6bT6I5W9
YR5WBqQv/dDBWrhtXoMzzf6ufaYcW/amZ0wy6ZIHwl8YkwMNcsWVPNDr9juib1Qlq7/RuEFD5HIN
lP9NNaxl+kzjcu5FV3sF5NNuYIFAgFn8udO0SYVWof0vsquNjJon2n3Deyj1XOS1uJQpvV3NNFSd
YdTT8fq0Q/Ls9pamySdOtHXTCm8WGib/lSqTa04c2msmIMn+QHpeURQrYH1fzz6li4iVI7qKKFIz
hZZY68ciWfpY87f0Xa51eH1uRVTTbvlUMSRlyWR4MjYifBIXKH4L2VDK3uh7X67N8Q6T9dfuUEC9
zHUtW9RFqD+onhUR7t5iebKlO9mUsrJQyTTG23gh/W53hJlMlxdGoXDQf5AF6Wue+5Mmyh1noDWj
HlcG9mY5s7qcaU4kdy9qOgKPzdGA7z3cS0SwPSLLPtsFP8ynGNOdTGyNsSwXOar1J/+khPSRQQrz
CmIhwOKUUuFB3swz3wp2+mikvlrw4bjs+S0UqCM3PwtRx0+yT6QIgHCuJ4r/PIRCtIca7IByLRm8
fJyVu5kXT/XRKP/PdfDk4bY5PxT+dApg5dwjlRByzkFBG8elBAVoB+cdMi7B/ac75qiknp2xcJry
yA7GZAn93JpPyhn7DxvIBXLx7qgtJ5ToLzzDLWNs5ie2Ua4nNhR0cWC3xzDnw9sRQ64rWJDeQ0lj
cvCrg5UHrXfGt5Ndy08mogOeAuMPk30XGfGMySNSVb0j/dUjobekU0FFLkHm4odejFQDj8EQnT0Z
9fcM36GnoV/mARY8FI+4HYFzPQH7w6QVsSqM9mMT5YLyabwrIALm15riTynzpOmq1ZZgQh/lNKVt
JH4LEjl8NkcXmGv/D1M723nLFfQrczq6QujemmjF5vUwyk7Gl0o9rdhUHsS+CFH4MAhU15fPRVbm
eDpx249EQcsLmUd9ANchGDCfS1xwBsC3WMxZTiiYi4BcuMnnFRAe/VxtTL0w35QMvl8rFb7qdjLE
NCpstyhM6395Ga1sS3GJH9PbEHLGmEGcTtwaBOzcyV0oe7CgHgd9n5mUE09CiD3VtyGs/ymg+lSG
wkoPraVCsVwuP+zn32R2+tHaAFf1pHkRhvuf/2vxNr5/M1xySUHmGlqe0G/pst9TdJrf7rS+apR6
Zh9iWjsOcdTBMEFKYWaA4qJnb8F7ZdpY5Jt5+clWXuGHnOq29Yj2GBTw2C3mpMZFPwS7s1D5EJLm
IFGxjdg15aftprMSO+cv9r6zMdb5WXqZDY/KaFo0h15cLnODbxk8DXq0dlwZKJyViacYxxeoDMqo
RDo8N235FkArlqJcQr0YHlXR9SdTSehYc7yaQPDguJCNhde8HUPJtlJgFD9T8C38fpb9i77DADkb
/0q50oE2QEQ45DABUhM9Vg7bexxl84Gs9ZwbgVc+JNqnn1hL3BhzVwrroVoc3APK8T3hSMmoECwB
8DM3yFACJXupZby34bhrnmkX5HPgm97L96vqsEyd04aZfhkladgsgWhlCpRlHe5kYuvartohv9gp
B99IQ5WtDlWBIYZ5lG5kLZOWgRAuqc8HHACCFebjM4YLtA0sVMOUvfqQ7KDyTeRAmFkEJzFFKo3m
7eFGNEUGVBwaKlVRDuUXbpo1quh4Hwa5TSxTHpxl8AbhKJfUQ4boGavgctMGxvvda2Hn5JkU2HXj
cKSbXzbsqaN2UkJZwv+LJh2kSFScmnLYgt9EIexkwyJq8ChojYpxauBV9X1R9z3g0jXBppiVNT+p
PayWScZR/XbMLeuA7eOI/kBAfbSTW0oWJU7qbNnK9+PtzjpOkhJyp49cr98BELaSnaOyPTkOi+CQ
vfz/izaenNmEiTo6533+WmOnQoI4q6X7b+kraZNuKU6hHVFyGi0ns5Ad62v6Gk7wwc26nBLR7ey8
PY/L32lwPrlpa7RqbtaQFXW9qYkHo+F7W5QhtII4bFFQOlyeAUniQCi7QnSnwVdbasGt7qC1Iz3s
fy12N0WSyDf4+8bevxnH1b/WJSknhAPjtgWij1SbErv2imuI+HFnigGQ2iybEghb+bsi4RRts8Ds
X8pVY+qXAAUXlnnh124QRvwL6yKX4aQAqN/Jmj8MfsIT6NltQ8+WBmAPmrJwNVsaNqIDKJ5jP4Ew
h7zDZ9v7V2nhKhtsmchOMGeBsunjHauL57+QISPQLDYSf/Psjx+Z4n/Bsz81vvetvQx5X5onGU27
JdPN6df03nbJv4IYYQ1z1Irz5/EkOn3N0kQKt4G2zM77kwS+6y+Pjau6kArcwIQ0PbAtlmYOVLXT
MmXgh/9n4+2YaGFIKNo3bpvyIz5L60SEp4mW6SVg4xyewIt9m8Q4RWaIja9mEHsXEtSy7g7ix53+
4TzSAAMLLxeD9hFBa/oFv711MPBvX5wrikFXQs67t/criD1ytu4/LUQ9PKeisFkn4Qyrg/Oyoaxv
2rwhQU6GOE9SnPPITu+reR54alBWIx73KOaJAnqNnRmq8DuVKS2n2Xk7AzKrrx0rLC+PPwvbdWps
i2SMBNgnRbVL1ofKZbshefAdlmz3Uf8UZ3YneBPiRepdkoghJj+QJZaaw4FQIGVvzCBpbEZCchV6
KNiMHeiryUpDOGWGgKPB4aSsH4w3MObV1M1iZgD9RtYZ7DGFbPZjzeNcPJjwmf+O9lVsOINTVlfE
ace9Fpf6ZcppJp8S6YuGGZ62RZLipJ/JHXm8tslttewTNpz6rz9w4Sgg56vCaesqZ8WvEh3JoG+z
I7nN7aWeT0yoTNKz+xmc2jR+3Juc9yFItgHbBhlZUdHYjOVwP/DBVIeH+aARlk82amdigagii/5f
NePTLN4Z7tPkesqB2if7ZJ5C0P8B2CjyheF+JHnVf+oxxDcuSKUs/Cs/ld2DfNWS7o10y4gIwj5g
4gzhehiZ3ujPYvev+BFh19tvl/abUlr3HOTrL5tmV8G0m4tsRACeuN712xLIDL1F3ysF/wYyaDW8
kLOnNKcM9r1dQmQdPPCErJ+uZkVZR2pw3OlE4ZhOiNKOrVQQNDuizllt6o+pybN6aNpNwlhtT9L4
vRjAQfXjCGyLDGw/530eSiFB34ysOZLUuz8rv4thHINxxfXe5xb1NlIRApPU36Zp0NP6izebVQm8
hb2tVz6o+3iaA7QLo+qV6tcHoq/LTgR7XmOn0ug9lgzE5xT0BOut4SWHWanNfNOhns2Em+l2ACcr
p7DOJuvkFO1+TaDEmEZVKCvn650bWpK2E1sNnHOE6ndrTWqwP39zL597MUAmC6cjJzJY3nLW0yu2
OZurXUanmTKEWBR+Txfg7oCyD2KIRu9MZDiUlmR8XS170sJKV7/+82RV6EUoC+8G35JFsXq/AmtQ
qVS1MBcnKGvqg470+92yYBhUekKLS7cytjyx2sG6l8yI8PyQyoLiYes5ly9Rox0m/0AhQkoIdokh
ywYoEbOjmPOa/z+yqnRi8ke8VqkUgf7/2Ii+X3E8y8nbYmQw6OCoORfVCmv4fQ5lvtAxv3m5pcYz
r27hbr+/NVmMbTB77n4TXHPyyrHzd4kq/8zIgdjiQtcBOqb07MK1mxc5difBsIfb4AxIcIIWVDl5
YO7LxPkQDFtgJUoDFIFjebsgo49lP9laV339o+wO70mAXw+7/2hE4IOJnFCtv8uF/xy2sv1nWt/Q
vxMTVtMK+HnSj+aWi+zx9Z1KJPE+mSNxrD3WrZ08eWi1ohKWyW0N/VQ3Hd2cG2WuHiN6JnW0d0Uk
O+IRtC9NDQRZ7MoeTiDKot2nyJN/jZdcpgFcECjBm4kaDyOmUjbVSE7Rw8tlDryqmKkEHHmnIJka
H4nortBVqgrL+OK009z2WXWlKpHDE1EXLPifIVtWPvqT+uvNQpbxgypEkGr8MgduMoa4/Ef9k+Bk
2GDbYnn8hC2hwJ0G3xBJVvjPdygw6K00Nop2fim8c2h8Z66xWvbTBfXeu9GVRVmRRli15wZCs+Vw
a9rTO4pfHJL5skqB6Om0Zv4E+efbvQHiZD/a5IIHTwA6e8sWq5Jn1McWRLHBDih1Fz1CVl3na3vt
C5aV2MeSNftI16S73oNJf+kY6kv80mX6D/B8q6I4LacAk7E4foFwXTjad9YkFIOErTmeWKzVXJVW
ioVA5OCJ35TC6kyThXL97VqLxyouCuVpGyyr+qLAKlVIYfE8Ex7yfBP91X1yG4oSIjMM25ObDyzu
ifH3PPnNiUEsEzw+tWCg6TqTxL4MV9u+yMs5XsFQEcorOe+lYZ/eYXRkLbk0wGyFBmIDk9IyEd9U
BnlrAlWTJLHfvtdjVZoL4R3p3lLjCdQkMAFatQs2N0w0fvC8nr4Rb5ZLuhsrlxEPdOqVZKdtcw3I
O1gHuDrCm7Q0LOgqbtolQEfCrUsXxc11FbdCs4yBxMt5j7sAouCxl0DmmRIvw5QGfp0+u0pCP4LD
80c4MdZwnWYmJU7E+8pYxR3ckbAjqARfEJJX6e9JuXZW5ClRLCkXYYK/amX9/z7uSz72N0VikGl5
FDhnZbFBAxFPlqTBI8RhmTc4rrci52Xj0xnTrutzAAl+d8HuoB4+JgCx4M9QBBZNamBxDsnelwY/
odTXIoBiQJ+YUBdBXNwGmWPItVr/jrZmFM3DoTSqc21BJCdo8FlTILighsXGXmYf+eck8Qw4ARZo
DRRFV5WDAzHJY0i2dsCRg4JTXgFM2bIRa96sPCUaOORAi3eL3gK8E5S2todYsdgVIR+edhsxrtyb
8sxd3qM65Rl3127wCrukWnqX/PCYtDbSpH9cIQWRGzU3TY41nVMmJ6dNTH0LceaQ6SRcuywckHVW
YUX79RU96OzE4OYofbBNnuYdM+h7kgPoB6KMkQrnNW1+wd0g8xrv2maFfeOq3g6/YIvHw6wvSNzk
nVr07CLs7pE/gEVD4TAOowUeDYenV63CqGEq6lONeIyeY0r55H9qTPD2bfoOY5HrMRt0EXX70z/L
B3f+QxeOz/3cmV5GGd5ddnFvLXGmWKg4OFLEem4J8b4hLX+zVdID2V/EMxfXvrT7WcZYfb6/eos7
tGcJ+w6O3wok9oNswQN0LXhQ8809a/XR8V2xIGrxVvZQXIWCo+qEsz1BgspCdpvJJ1uP0Uvvtkuy
vq9pXnrZ5LZfTsD5cR5kkDOiDYw9PuyZ8IwZtthWe4yn/HtGgMzIfAh2ZRDzdmOl5fzufXA7B1Hq
6Lz2O/HcQzo7RrHpXg0ZQfoBeTynsSDlwZ7L5PlpnHxQf5QmFHhSb5Wytx2szH5PDQaBx0AIJRBV
bTFn28lvIR8YZJfOB7HYRm677RxC5iVC/GbHHDKbiwea3h5S+iSRfjkLIukJ9f8ds1hLpJEkSJH3
b1JY3+TPLpDAyVcJEKWHaRv6kz4jPaKOJhZzhLJVxWCz00OQ4Km353njgdVAqGmm02DYy8IQvAJr
ZcLjRPSQ/Ar15CgKum7pNET7PAgUVjggrX9tkiC1Ir/bR5rSJe/hIzwahDi0SfCqSdeJroQBT4Ez
xIY7TUBciaJ7ML1TzlInGEFwd4QOlkf8OFzjoKrcNDTwe6w9GpDfLTCJVQQPorkjYE7b7dwdu23E
wr6pTpzlKez1Aj6go7L438ubnZ8ktpjYj/ONHYaj8cLBWhq7COawkZfVJ4rk19HI0x9XtHf2Rmqk
NxDsEfkm6KEFrbAqrko8Im2+wigwTXXkPnYW9jIo5LMjqfkSzlDeW4B1qMYIxxhCDrBmJVurgVZd
rf27cD00ZAvPycoucu71rgI/UpeTpDknogohZ3Wt3L+VjSiN2jt8byKnQVgA7pyXpNbTav8gJrqE
eR+DsYH+vMqBzMARISY2yq0MEndkPUXjUQSu8dj1lnoEf4Dod5NOCgApgrFjn96GOFddcPsMlv65
P8m2vIJuHR2fJtxgHjPCBqKyMhqYY/z6ScRr5J3UjELV4mkMQBN0t1rdyVzgbchf6I0QKtmYJkT0
o1WfZTQi7/fD6sajwFuJzvHpdTnNEcEzlJr5IGAXiP7reUl/rpvqCemioE/SQtceRiKKZxKPyH/w
P1ravB542uyrBq3oiMev1tu/q5K+b1GsDvB9IkpTrqztILKPtELuQiUFKQyHVTb/zomw7ui4r6Ih
EIobOYiwgVUBZcN5Lu4LUTjmq12wddZ6Tuz5s+SA0CzEA4LfLkEygaZ5LbA0rHR5INvRdsKLyUTT
RlXqW+53OxVUbk9lV5+s4ePLpUyJOnL31shneZ4LTr5b5O9VMzB6rO3eDQCfrhdgJl69O62I/2QC
qu1k9LGUPGtuvj+NKWBZ3hwYyGjMw5JdLuyLqvw+HEFV0Ap3li0bmz9bc8YMQJKXRfETcxjzCe1s
0/tjYKddDQRFLDT6+DXJAPU3GBqWX4hkdHU5glykQ5/y6NNaUmeQdqzfOj0TAwNTXzRpHGS6jS8W
zKzWWKkEMwbYV90V0ErTxxCSqRILN6OE0VgsJwxQzMv4WvMLnsL7LvadEBFq7LzH1swQoJtUgJI8
5WB5rPmWQ3YnLqZMWNFXk5b3b99W1hK8f1UKCXVBfUbsG087o4fMB7Ps5KHaXbCTYbOoB0E3lkRV
hWnq+t1TGo2CUtU+IiOoeACzeX1S50aKyoLUsl33jKsk/G3pqWSKasUW6lBMPXB/wyqNEauq6hoM
tGLEbwXfwo7m6C1Y8ft9xGxyXkItKXfuTrqDsV3Py6nbxCtJLEX5XF3qPikZihxclSZa/1S/7axf
0MYTrj6kd8so+sZ8A0EwVqr/H92OJLM1dsUdtFTpRA3CtzHFOK6TgkWv5wuyAEsSO327TjM/IlBy
SkpYYHG+ZQ5o5rG8riPTBqv+PEh3C205mmkO8xnV+XzdJNkj1wKxai9q+t2l8zqs8aW+wxRQClyV
ZA1JoKzM6M1kw8XOYBIf8bEoUSjN0OVYN3IQtC7tSN8U1pxMgMS2p5DXyv0S3SHOL4AyJmXcVvDK
opnDm/P6PL5OFyb8DOvaVPj6AL+eG+mqJGEVXM8CIN5W31GcvnUgJfko/9XBVKhcOeiJGkbGQ4lm
Wup6lugojbrIp01+KD5MMmXkDn4WieqZk+0VKYs/cBmblrI9dWdrDrHeTTRQe1tVUGUwk5ar9YTE
cW283Wle+xkkz4olUp6TrFkk3mE8vVlXrRSIhIL+OqZImNg1cZcVHdEj0nQyKBRhYlY+PingHqe6
VV0J4S0YqgE/J8gVn7BjkWmqQmfIQz8fgwFEg8nHlILN3vyJBYocUPag9VfB7QHxYs9H9yGQ8Kst
vhNVyQSfb0/wRbGaocYT255xW4PxwjOYLfgU7xgjIU/WFPeU7wc23tblbn6C4rT0AWiWKOa/7U4E
CkcyO/iI8zE9Y4CmesQcTo6YCl+LIj9nqkMeIatY7DaLVHWCdAMc3tx5YQenwO7rwfadHbh00rUX
sEYc3VavPp/ZsZveTyOTQuGrLU9t3qr63AwwaFA1QybAkp59xCFop86WARVcFNMyp2oZlfFs4c/e
Q9Hq7rUuPI84kUQLnpk/vEvyHoQeH6soLA6AL8sv2DMPja3dja/knWaRIjeqdL8Sbes8QVf9gSmQ
4RfkdZmzp6SiPkaQkW1VfSAqwK80S4DXVfzOXCl5YEQTWxFkuTpCnEL+0yLFdOvn8wrsOdcVGJB4
HC5v1AxDaLt7Q2hsKonK5onrXzj55clmNIjgkm7+AQ3UVIAUdqqEWL7vCVXs51bivIiPrCO+mDg6
ryXHuQQ7kbAobi+WMWGpp3bcNUDfL2xC67mAQoG8AOL1+tWYjoRU60PGx3hd6q0tiZ6Nin7gS/dM
EFZiVDqX2EOOtBjg/7/f4kta84Y6W7RByjSP93OWRH1PhGcAgwVNSbTHis96JgsLGBbhYMMny5zS
2Tn7HElQViEjOOtwgkSCpRywYI1Uoj0AXBmTCztwPUKrMS6oKmS+SY97yRPxOGl41PJiGWD8sJRC
T86XBtWu4JGDkyyNMA6F1dar7RGiIOfTUAnKx0JJug4qtu1zb1YSCnhJuRcAuPuEIAnuPJQ69iD5
ylm5k/++HR3K38KzUehIQWMTWUHYGmkAoK58c3+qW+FcXwjrQMoPWwqmGCS8P1i2X5fTvDcWdG5U
U1g9g6ANLCLCsfqGJCzIbmmIpTaOFTQajN1phC80KJ7fTduvpcBE8wRgkOHveqIJmCK2FawrigwU
oHwthejcdGtK4N08Ica9uDR8D6gYNtxn1+jZXNNgdNf+YMfPrIckm1ZbXQL8Xf5Aq0Wct5cCZLcn
suoMlkYFLMBAEhGkI3ddri6ZlyPwuj8yvOw0bIhU4ma06hMb2g477GQSwb/IPuFjsPUxBkUSP1D/
wmkEalS4hEOTIutq6D05Cj0kJEXfdrQvZX7KclbGx+Qm8pwe4QzL5057QTDqpbpsnEZ5oDwLGr5B
PBFyk9xgx8dw1CaZL5HBpLwf0CNy+/9c7Jyp97h09nkeb9HEhdmzXM/0q0HkpgetYTDFdGGvXVSg
VKfBlYi7bUfINgCLbHO+8vfrHCQv22crFOLnoBp0SPrZXl/0Ta9BogcJnDvVFsBk6Xt1q9iWDVss
yHdsA8CpJKKm5Mn49rB2S+n43XvqBTfIEO/2ivYfmlZz09clJGvu/2dUiXgCbkz0hcfEr+zREtU8
ffwC0HOJ70oOfZI7VUffPzlV3Akq5IV09HKMDtQ4B5aZwBn7dMs/+6wjMphTYhIpC2SczMKFkin1
vdEcuedT6+BYvQW6bGU9W8QWnvuHVTS7xtFG6Fv0LrDVRobvFJC+iXkfZ7aafyr6ZsyHO6eqE/TN
S+oFgJbR6Kl3FwgrUWtl5J5l6GErhRy4pPCUJeUvXBikcZywZOVAMGxbE+Cz4bL0A2U+yd8NjXFZ
G3cQDr8+mTwMa/URuMjS/F5NgKsUDkT9yaizHDCFplIv1s76LmAbbwwdLHsEw70CFGBPwsw+nnh7
/qPA1Aizqhc8vxTtczFk4wgT76jYJlE1+o9GsOiWDnx6qB75n7bP9N3xeg77uugQKautD0rCky2P
W2SapdbqEAVJzonx/SDe6ilJZWHZXFF2cAZZPc09aSWG/f7mA4skE6GRdoe/rcThVlFvSJWuqfuH
BvPMhq5JBCHC9Q9yMnEA/3Oj1g8m58fdcoINeB0NdEysgl4J1uMKJkbCiEw2GcCm8/m1vN1hAy/i
b2NQkAc3yYRTZw6nJxq6qtCdDD3BBEN3k6UUTu7ysYvDoOtieU6SKwN3jA/GQFiayyz/qToLO5J4
Y3r0q8Ehs2u22c9Kqic8pt8oZtqRZG7MNWjC+MT+Vo4PQfoaa4g2gKWk6iZQFfY/5VuDEuK3LsQI
iveX9QLiP7WiEGpVKe34NVPrCXpGYm8V92tkmJt4ezeWk9d7IiDWulmGUaPgL7ppR/b6Osr1GTr1
wK2YToMTwKdVQkseFOTUuJaHZZP9/+j2VXy7Y2pF4+T7p0HvF2qJv86qu3WE5SlgNehgu4TjMDVM
J1fYtY8rM3i4vOTzLkuuPTs2CmMjNg8IeZeR7CDF8xFcQjJ2RfNXiAw9Tt/yYzALcH0GLzu3rM/R
OTFUvKSyj8Q4muUWOwiyRk2sOqnsECvZRyOWbYFMm4eaEjqRV2liWzhdu3wUC4I29QGcw7ByUZI2
Pi05mSWoBQLov1q+zOW3gLO4YGyEJOyiT/u70Ie3aAGEr+BaFfKC2WmzgMyOGliSwUynKaWgxTBj
HJsUbaJnb0j3x2M9iQs7g4aADitd9j56grfb2fL4KOi19Z5vYqciJTDkEvbwqfWByuCRcJ2We0wR
bwTjI5S6YHB2r3uUv47gmQS+iWN5AqEIcmMpHpNt9JUI+pU+RFKkU95CLKwWIyozvhH+Vh/jRwc9
/+Vfjrn59RH3LXUlr/vKiErrpVzTsRKpupc1CO6ZoALI6nilvQQKdk4qvc4KzReEVqvR10xnLGMf
YuEGdmy3YE4yuaY6VfDZ8SqpQDdTg5Uzu+ECkTt5dbU8HQEj1lR2SdthUfkctG6A/Io4+3ohNm4Z
qKV7UBDRg0evq+afeCWcb0xwQnQk6M2Lg6793CEt9Ru3zcX9lWZaFYVsrVQUBY9NmAvd/CGFKTD+
LPo81u1itajbRCSmJOyiklIEjJSC3Y6Ljpd2xD9nJMJGo4/ynl9zSnxPCVZaYbr3scYQ13oKVh8i
jpm044WEukh6k9JLm7HjdYWNx64ThWtQK1oor5wNvwIRXN/nT5yR0tV937wzR74wRaZgjjmb/qS+
lxKV6Ai7HIEs/CYep3vPsdi67ddTDL1vgICLrx0vWETbjZItdd+8JMvUHah5mBB/CvuAnRDSRkHd
Kko1Ng4jId6NgKoNedIcSpz5sUtIiIZdEUV4NpITuyn+UtHbzgAh/3VbTXhvsynfBlAMJdDD/ATa
tsiBTfBoKg0/sDEKcWXd0gbyCsM+M4DYnK/FInvvLWZoUQYJxsS/MMegYKOWwivh6TT4W/oplRlT
UGgWIx2xDbcYuS6ll3+4gjLcmRRYf8CLHI5xaC8POxmLydLvG86fxcnRtvWodrX31ZTo2C3qkso3
HbHunqVTdhu5x24T2tR//8rNFcS0QvgYLSmJbh/FyvbnaSlNC8f5u7TiA5uGLDbiUMcokhWFkHcn
2tcDptyu914XHdDQJSZVAFhIBiILvoGSmnuj1udf0uQ18Dc6EQopEv/md2xsGavW9YQ0v7n4DqXq
yxBpu8h5peZ3CzdhvFQKRLcChEvnTeKk9KQ+2GwQsQLX1KkvmSCF1W8QNLo23EdlzGyyV5kXvm6o
ZCKv6kpO9FnfpbLIp73MgCvH6X2cUWZI1vLhJKQBAlF7iHHfE3v87cqgj8k72DPo6Fxi2p1pni/t
GZ6Gs93oGOwcikKakDPbkOYBPIVX1LVphySbEOcX43uUfZ3YbApWkOShMn7jfNkIqU9OiawQo2Un
XYMpF/TEDpnbDaQg0suKW3de1FsQjbjwCd0utLIOuizq8VBNgPnbUWauaPrqzR7/rt+cj5LSDqf5
5NuxC/elxnaPywhEK32Sto06dRVpVM0VgvZdknUFcE0ztAc4HvudAXkn3lA3Gwul741ClWQ6vpOs
QkSxV+EVgf2vctAS1CUH2g+FOhIkc4b/sGvWQNv4bmWPi6CcG7iNAH9eTEU8p0MGH2BF9bLTbQrf
folxTHTgJx3Otb3V55AUBCvScNv9wrfOYADKF6RtQHpMV8EnhMs8lHUprxafD8AgmFRdmqhdeCD+
o+esuajrf6aCcYhtPhHnYLnHT7yCIQrT/72xPcUvBz+C/h4cOKTtPIJDIX/8JwfdEBRRb0vRyK+h
JHssFOLF5cVl7OPRsQOJl174hXThDOCTwhZWccr5PoRHXrLmlUpL5z7CF7BpJ7d/xMe2kbWBw4vw
RTBMVyWdASTUOerZ4Dluqoq4n4Wee6U2JN24hUfa0goQPJs6/Ctc4B9Fcn7D5cGBE2NxCfFIL9lu
YadycEs/0kKXsjphZtd1WIKYSz3ilc43I8FLVk69mzRXk0FqWGYb9l6H3zEbNCZZzdESAlAhRxWr
P9l1/HtGLXLP4/y8ovM9+KVehzbEGGeWAcUa6RkCgPkWVivRPI1Te+RBjkThy8uvjttWpaYi2Wf0
GqX5u2Vyybs1zfSef4ZuE+sdU5xI1QwJClPz3BGiYc8W02I/7Ny8knZ2K4iklCgccJ8I9ytttpHo
v6cVBcJ23hYt15jNRou7qVpAE3WjF3IHfDENqB544bV7/sO6SppfviuHTJAUtQ3OzHLBBHZ9tTzR
EF5UqbOGQfLTRfVNkO6WNbOIz65ctsf+4UcAI9EjlqSTKSGnWClHV3H6HVAvFZvJZvJuyDU9EC8K
g8SERiblevZYQgwaBN/jIRsUd8q488U5jwEPxfLKXQb3BCOGEzBsDEOWQKGolTu9Ya8Um1ypHtPx
mPwFBKd+VdDOUIKiy10H4/ajo+Ac/tuIaeHiTWlVsbk8psfITaBDVPxCCAC1EO8FzxJYsOeg20Gf
hATgli8dsmeuetsoj9SvHNJoPgfu4OClkx4CsSzwR0CjUat24dkdGrFv7ANbApFzRaPfyiILY8to
OBSbjOpXh8TyyKVIzjFt3gCphTmsLV8SqSyMmATL/M8rJL2sHykLUa1yO4gICDaLEmZAUUxnHRwN
bD/LgF1o9g4OzbcQwELz1clYFdETm91p14OXUmlGbYsK1mdnF1NGGpmHGISasy/0f124U9L7/5ZT
QFrd/EzApwh/ALpEMD1Xng/JHPWwspX3EiADmxwY4APgocb8y0kEc6MDV7vSY4x1r9w+S+RWqJQ6
14Hxn1oOLS9WDKQ9Qk8hXLWlvW8go+tmMhrYP230+XZcyQByNAfL/09VQU7+DpirbKXNGq4c44pF
c5ch1DV9TY1Br3OsI6X99Q9yOwCG5xpvf03HpbhmFi6yJsSq85P1zbdOlUsgD0qtERUTttit5TXn
C8vDruEZiBTgFlRNuTSr+7mW4JyNK4FAJWzm+5SzrXSyuog3zJ3Uc6N6cKlB5XLPA6LJ/MFE263v
pNTMLk25kM7Id6yqpjDjdkkhNFQaaiHd126QKrsj39ufoPgE52MpE3KK4Izh0sEAmxkmoiusHZqV
6yJ3pOwJox0uhDebOWxoC5GI4CyWHJrof7pzA1GT92NyrqlGL5E1sRvLs61GSCHx+sgmfkpDurE+
Sqn4sdXjxVkMGLrUxjO/2pBBLRDt9BcCwK3Xt5DM8wyl/dAxlA4faK0N5Croh4wjbqpjWCFPd32Y
7itI7w9/gZ63STZHTG2imsJ5efh3VxJ/f5quWV+uf0iIFm+O9KxRq+SI/quKecsRkORhUJHuOPa5
DF/5aF59Je/+WsulnOoz9cxRrom4diHzquhZIY+yKSR3DtJq+wjSlrZ9Q/APF5IcE9fdq4JhNB3n
Lg4OaMngAN8ic1LEiMngndIBFgWFfXGw/cCX/xzL+PjaLcKlYWFZB8QVT5KQjdI1TpKeslj8Evqk
8kA9dSiObLTkI0lPyb4z+46wUxISMtgBJRAScJ0kaoz6i6xYhOhsJ5JRrPuhdeU36Xx1RVjuG8KL
1auZomoTncpq9/V+/kvA1OjU1p5Q35kHkoZMoKHVQovu0EHlHE4LCeZXMQe+a+KofTsqBUrdbscD
M1jjIgJpNLUfUiuTirpkd8waGoaKyreNQSKAiTw5cH2ZtBd7qQiR06BPtuAHyt6KfL3j5Rv0+SfY
fxeIn0/DqNBhHwYkmfIZe06eJizdksXirHHoAbeJq4FL6BWiLRaTOe1IBFhfsnhwR/Yu70gMKtfu
oW23JEJfgNygYfsx8AQgdWKejiv4L6vt/31Zo33J0hOrUr2fyZvjZyVG6hUiFhBBhxn3LpwK3N9W
s/ogW2k/llpoXIhGsokH/ebgIHY7olb35pVTzEqjWOsLSST9Z5cHQVo0jDbd4J36wn7gVKJ+y6BH
gQsUkT8gzw9oNeCNB2t78KKcoUxM3QcAzf7nGsFli1OspDi6CYUgGnIOGRJPkNTP0TIZFUrYqm8h
zcANFNey0K+fNPoFBoYiKuDqrIFwqhBDMoK1j+pq1yhv02Jv3aZUoXwx5+lcjSTuP1LhraG0eiYe
/9DXfTaqgQBMyuwC+HAz+VGvjfw/Plbj5WqyauB8QHDjbFvIy5A4A/G+LcNCSAjc/z4NK1R9gH4X
07eCBby4Fb1QxKIQsLwD97ItSI8KcvTtNnWc2gAO0fRsEjV/0K2SMkEtgsIdb5wSWhv8XfdZF9uv
MjaRIdD7YkrxdtRbmlW7DMm5Cs5+HJCsBLbGNyTNRBaYCc/nPAf8XDu0lT8L5d1UpZouX1wgcvTZ
UFXwMX0xarpVsJpmLIFfZE9eForkAFgtPYwVfI7EZx2tFP5TWzq093Lo+aym3rGS4yvLSnXfJ3f1
0roV0SQTCzEdoXLymxLmNtmDwz3+gVmY3Ju4vLULEGrYtSkwyAwfHfGPPiWubx7RdlCXjv6UdlY0
FlHxsdPUysQMzliKscIAxAvwVjtFmPQ39h2EbxbQDHRWxa8HAzTzboqoE/UoXlYShelLsnnwySMk
OsNWbG38L0vh0VuIi2RItsFT5miRwNLZROQNUVpeXNJP9v8Tf5dH49cH+uw0BZZHDDzcPACV8bwb
T/oURWiD9bzZo8WXer66NpMeERKU4ujAWTQqfFcIGcx2taP45O6Gll7eJlwMjoNz7hv7n9ZlDGSZ
YxPp5QL8RsJBbcGnDSDXb+pjUGmQel3tEMlDSwCAyhQd+dORTefXwSV8iY4cloKAwfWmk3rvxS7U
+bkPRd8QFYu/RhA6KSf2CUbwQvQdRQpuwx8i7R6eI15TNBxtEkZv/oOb2miHJDAS4q6LRJp5EfkB
aFXEZytrq+fo64J11V6zAfQHywqDGpCCAsU60Y4hLDODiRH2u7mPQjalEfuP21bonEE4veVTAjUM
76p+iLJsaflx6bdLRDzC1UmqoPlJij7iOF0KuqzCy8cvJHQpJTiQtJ21seePpJg/yL1UYLp3lEnm
xQwmiUfrIge2CPrx0uUEzNILUZtlTAoMSYZoA88M5Rds0bR8OBTkvVZ5P2rMpipYIEoEYQcC8bO6
oiYfQCvbvnCfLxBff/rAf4Bdt9kQ7DfjQLHcK7/vBKhZCbEG6+2UbgDBmbEs4hPVqhgJC4FyjFwx
dUzzDFTxCmXBNLLz0iNqTwkjvS3K6VepNFY0dz25h4YFXQiKY+PnIRG4bXiD1NGeTX8l+GUNZZmC
pTHwOKK35esAhbFiF81fBUM1KxMA+GofcPGaBemXaURsj9Qk/QD7HSdD7O8tpKfADXybf8e2Ei6Q
3swct5k7Pgk3hxByme6CI6L01twFDP0lvtS+54g5jJCSx0PqJPUEYwP9hHKhNtk0Vtkhmeg5RRwf
D2VgwWL+9RuadNwdlyceGXzZ+MLXdbRzcuw1abzVoQZGp69aslNO2jpkMqQfzPuvoOhVSZWuwvtT
8zHeDBNYYvdCo8qLGHyeYduzAAQH76iOsv3H0kvxnKSbKEkaYvwKcGgIO+Lc2d1nPhc/9AJG9r+q
hBznRYhLgHHaDWhuO2ysIhZLCz8ZCg3793quiRAKbDT15qjHoStytRZglPW9VZsqWSnCpy9bcLXq
v0NAq17yL7qlqSof0xN1qlq0FsO1Lr8+VX2aUpU/OlDz1FV3RVay/NgVNVG9x5c0QWSBbdePuVpC
NekSZZHIpxZqaenE4MsizBYCGBPpJZooVd2QMnYewa09b76Op033PHNC0FSs/ebCR23AH3VKPGyA
bQ5SzuNcUY3v0rVP4MAAZHCZPXCGecnaJ4Sj/vZlh4hkqVZHH891mSUfPJeiQx7SNg67w3qfF7Od
v5RwO78qtOF53GlJa4bUBj+QHWlqHcwVY7CmVCYP0ToumwAgo25bHlEYQKKHDinYovaZ/faoA81a
97Pl9XjJjW9wndJ8EMdw++VR/ebfxjkTiRbJxuGbiL7KfSLHFBh2gLbroCD+aRtZPwtCqJwDs5LI
PvVyM8MA7qjl0RnRbIVGouT5oAWp3nqduxRShgbcKjif3c6XWFg4SacWw6hkLc85zJ/KS4Aq0MB0
nhLJVyLjRbjINdZwNeZ6yAKpMJq7N5jajuPQGQY9RAjSAOIkmWGNrjIxCCRg360e5YFsNxAnP5VI
8ybAyTMILhMcfACI8bISzu13QufMhpQKzFH1820ElE9h4kl6ZaB8E2pmTh/j6vlghT3ptQuD4ZhT
YfsBiGTwctHYryfzgwsOof1O0s8txPv6RgMia6JMb5XK0HGA0tS5v1LYVz3BXxIW0AM6R6aXUaQN
mPvRcbd1xwCWvmQidMgtsDmZB/L9ibdy+YxT43lU9Ll2HkXBYnBSFxyGYbfl/R+CFGlj3MvNO0rd
ZLULB8jaRPyOaJrDPxlFXXFhvy/97Z0Tg2FxRBxMz/3k+2JibMcm5u7jgwZtPP7xSzNHJ3gYo0VR
N2yT38t2l+rb0Ew+myd4+r636gMC39lQZnrXndg6ENWFAmI+B9Uub6KtMIRUJTGh6YZMyMuPq/Kz
Wy1VyAc5lkhTbeKUDY5z8O9scCs/WibqLn7yBqb8IIUNPjGK3wI2PQbLvRr1tpWXZ3N2rG8F59d2
YqKwxmirfoTmRZidYiEP9pT3+a2lodMopb3XrUNmNEzZsrkxqDR2gyC7SqK3V1j9/AWNxXgbsum4
fq2XY24KQvjgP4O+gfXwPeIZgwr7OohubUT5Nj5sQR64Nk26gF48WEV6bpT3vb0ETntuGti8/atO
zxBruf/KUP4p/uADFFZHBnBMzY6myV/GZ+ixOWebiFnN2OK6g8R0werXdoC/cSYaKtzS8J4+4T4e
24WsQsCoM5FgA8Ub5EjriNj2jXGbFf6Z2vM+mGz7RHoMVp2xIadHcnle6oWYiHKDQ/arLSaKcfRb
DEG3Ib/t9aN7yEMwJki4L20t3bPAvSaiUezvT8Egpb6TF8ugGJLO7uN075dSHeLYcBqVJuexInqB
MAYXlWBGN7Cu/AWIH48t3I4pBwg5LhZSI+YpnfQl2jdaTLIPxf/5Ey3NTnP3mW7+aP4f9zIeCiCW
7avyvdLary8SVcu7H5NNwlan0SzM0axl+aNbTv3Y1ckfwQ/0K7b+Kq870hARoZzXJ6+vBf1dGWVz
xluT4QgR5CUEXA4s8QRBSkL82GNIxVhvPqGRNeQWAx3WWxa3lYuvBPuHjxpoApuZvpiKmTqZw6KR
jRsmWD8ouejSNND3xAkU7UgYWcaSOLxrZ3vzSAQRedFEjvvgpjeGmZ9W4HVYUSkEyLLn9IV0uXvT
BzTQPAgNY4wp40ZIrdOKTRqyekUWeqVfuggThpf4Bwd9+XX9UvDNUZRn/qvxl0oXjXcOpH45YcRl
wm76nMPaQZG1fDCZ2GXckYZpoIE10Fcg8GwNzxcWZjckaxeS/hVQhit7i5/sF7d0M8r8KuiT1dG6
qhlbinlmJh7VV/d+q+1wXGVdPCcWIRqkVDMAeEX8AteHIMjWCCbNagmcylmOaWm0AwN0gS0tqfgJ
wGXNmDwUefokfrrLPYbCTpAkpSHlmxIqL24amblMx7hfiJGC15xDAFHc8GmqRhAhHCWUIRWOYWAl
lfR6dvN62UCSzJSbj80RDzI1iwjlNCGQd41ym/ColQmkESyCGVfgqCWRJ33uFoRfHkrvDuetp2GV
5mDaEO3wc3La5QgyGnI/PRtmdgemKmYlF47ArLR7zUrdrno3c4AWNP2MX+gliMcj2wsh2f/VdYtQ
TIK6VHfsZph66mBpoMrzVTDRl42v1eLCw8tHnjtTSFysAL/vvHC35V5+itofO+YcXe2qYHGZS+ao
1qi73F7+5wTzaVAG3yOVmTjrQ+p7jcLMd9EIPOMOkBvkyHg5HRafTXtBfSyi5U6ZPMxdC35qbJzE
ooliaMkwAPpE6ytVnBmjy5YeMk+YYnaGZ6Fcoz/1Cvi35s3iJrwvHdxCXkv7g4FEc4w7BacoN7gl
Xf/nAbmVxfBvnlDvlIWNmIQCepHxTlZukPzfhAxcvA+hCWFZfQBQ9J1F+VrcPbgcGAB8968ubltM
DJ8B60FSFM5+gEVDQ9pk0SbL+BnV0u6tJcM6BmVbM9GUQfR4CE3TFUveAtxGBFesceVDBNukuBsQ
qhbksFUCPUBEqMd2eX38A5bZAWvch9ntTlRpwH4oP7R97LHvTt8EIpDA0rAWPJHngqMw8c7IGL46
ZfU76qEgYSO+Oq3wBMkks5okmVYaQsI7suiHXgSxLkGmmAQpdKwci0EOe+VMLWJ0DM8CW+KqjXAM
CrIWS01g7m6ufkhmF6ZrDsOVZN5UYk1PYz/Jx5Rw5wHzQ/bxkIVzzcdqvNdASphOUEwtoRa+bY6M
aQr5xwg8YaGo/vKyzbOb8u/mJ0NTPum445HkzrJgYQOGnKCWhsjYHH+X06NQLdX8nzDh4EodV+sc
wxeX/6AUrtyGqR98GXYQVyXyhZQ2tqWPaciSx4yJ3+DvEDhBMgJBkp9o0NYdmbK/HoLcb2HSovLr
xlqFkDGTLPZONZSy2gdVTfEmieeq0f3QfT6XH522iVXO7bqSQY9axz/vaRu3rvq+h2Eik6QzxbGD
4L4d733cUE9lRFRQSg+m4oIAKWG7nUUvNchjElGfKibul5L/v/Nanpn9BCbHMhzFZBO6ZE/s0ByT
Lg3bL+pCx8y2XuI6cn/s5WYt2ChwUAsJJziZD3GAsEbNO4k3/EXev7FOprF12ZaY05VSuxQ4Bfif
oCN8/pW+W74ejeUmbSA/3SDuTS7Hn2lv3dzURw7to8Ln6BBL+0EKBT5X2QWttCX+4AXITBFepcsn
h3WPgHHek1V0iHXmp1LS0XjxN9q43UZ8C67QQgXvnJpCuyMGYr/3/eXW16vpVucdrtd+sr31nP+s
8qJrC0yXCequET1Pk3oDLrtB6zKZlR52CUKANwpQvFlaqXvZXe/7ISmxQfajPYh+lO/niwei1AQY
3qRrDfE9qyaKJeNNtZfxAuo5AibG2Cu4gOIypI4z3UfGByeAh/nvRr10W4+vaw12nVEctKjLMAZL
7ZgW+KscmTbk44AApGcpGXtsltwgqzxh2u1f6zle3a8e98T4mzMU4MAscNcwvEAtTPZWbLdB0CFS
rbDNFBicS5C2SSWGlxNRHjGEU8911CW79JAXaWUtft7Z2i74EGWR7PKDwMWnxE4FUmkeO8FaiVfn
u7KKF80iaOBzZnZgW5ElquUcPjh8satg6pYwkyYyX7RKAv/XWbf/8xupR9id0g2/XuXZjZX5qf0R
erYv33ioslpala2T3S8Tgm5sGfvJJQsexfU8dMof/4pe0FJtuSLSnco5DYFgEFLt2pkB9OhrODEP
1DUR0+OQiAK7N9hTGgrHI2fsTZEEa3wBuXD7T2THLI5CojeosdlTphwhdhTUcVnD5tcXZYI0nQJ8
NQ61SVbopdecQb/NVxJ9xLfc28VvdMuxn0dJH3adI08bs34Q0WZyFTbKC4OgJVV1KI70qoH/Hsg6
Z35flD0sVpi0JVl3+JPEMQscgp5PU5svmifMfYZKR004TluAfKbC4ja9tfmrMBQ4zZh3BMpz0a4Q
O+QPzRb+NQ3uLClWcx+m2OvG4EbUAMf+GLqInpef3dFkwPx6O8SDSY2rE6i8baisOKUXSuW6MP15
tNnbYuPKa5w4IrbYrbPCqpukep338j3dT/K4VsOWB134vQL+w7zEOd+7W7zsjTcVnecsa729UtqY
SKgLiDbdQCGY7NNLxpQ1pczef6p643J6bdzDvY8DKij+PFqvI0zz1d0U4wdZPCQpzvM+aq/DGS3y
wWMLXXGui5VBmvEF4OJDA4XbiAhO+wNT6qDaSP26nPSLI6VoeAmKcta00iEJvxU/irdmYrksz1w/
YjCgxFQvuSLl5qIZCU6f3ocMZl9H0lpoDkPFd7qrvBFWf/OfApUb556dKMWwynbn5XtBv4Ju+8uR
Gex+CJmp1h9RY7itl3Ix4+zbWO+Vq4PFlWJpIkIK0hlBE1fQrVflOGW94tk1tXU4IcNP63Q8Zvzd
SnxMRMConZSCHQRfVAmT8aT4+J6Xlu+jDU/YoCXlsCmS63chrasmT7yn36XSbJHa1ZMqPjjUA59H
NgAIwzWSlwh333+B1KW1o0M8zYPRv9qWPgdpa+q6Kr1/gbjL3784lXp2duhYejtd3Ts8EKl7VMLe
zyv4N5ULeBWa0aDpmWDPS/NyHrib62iPlcpnKtGGPkrjWgFSHG1KvI0iddPnFxaQFg90nf01kGqe
J9VGbFJ304VSLrByjiMoIkcxwb4sV8AErxdKZkGDBDTE1PM7/aRPiUw5t5ZE7ooET1iYT16Qf2iK
e3QOIV/1MYPJh1sc8ndSQx0PMhb4PVwIf6f1Ycs1xu31jO0hFlwUoc4jiX2vI3gU3+JygjK6sIhV
dEMWZcvnaYkfx/cLvWinROjBmvtIz+l39Z98lDE9DrAwv9fkQg/zdjBtNi8AyxuX8VCZa+C1YysT
PQ3Gckt7V047YYM9cpCi80vLG7eOh3z9DwLpZqo6FxPSIhUNBc+TEWcTP+XgKe5lrX27atHyn89L
YlKIAI2S3CKAeWdarjDH+gSLUYk9BLgKf1P3KAJbCO8bvhjDDMg8oHPGiH2W7YeFfkfkIAcB5KBa
Nm3tW73qKV5rnKOW6vlfXa3ljrb4Orp8cRj7jOXhF9oq1fAXo5hQbKJ2W/Ptc42P6rjYE490xGm+
16zf1WylQtGE9f1mnwwuD7CUqiNLhC60RFGYlk2VKXRQ9lc8BYZbJ0PbQxSpsPJvna20Lir7/WDO
iAiDmHse+Et7TSw4+ylsxfzZLONbxG3TxbrTfXnlvYyviaf/Zt/KnxnyJiO/1JiymirFG/6DV11G
SAF3U0Us9JJQPTg9xWIRtLFLIH51Nrb/EVFQPj58q2UeW/Bi0leTakxRnY7uuoLsndqPAWQbWILz
S9Ewo/Ieyk4tDmgF046lq6cXbf27NyY4W2QoaiTw92s6eLdboIUEyieGhsCMqvTz2bFcIuDIKySG
iEvPQ/qCDNC1p1DxlEw7FKVioQCQPtEm9dKJDJ9ydH4PAHIIKYmkTTaZp+27AXDLhmLi2Fp30JEM
PPgNYbupd17DKbT+z2mM2nB5JsTIX7x+sEda35zTYefmUVaPTawz62vgTyzFC9YVlrLWh7ECuveC
Ip2bqV7DRUoVAlCjdWWPdsCN6INS3szjeG5zrbLOf3OyjldkK0y8DgXhWKW/yPYn7DIpnJaQZ7eb
XIILXm3WKBu6NaofdmeD3nelMA+OTWaiOjLWpnUxyE8lvNhnfPd08Y4AYOnXcScRqeZsHa4rIHPm
uk/uoq7MDbRI9WXM+uL9XmllvPNBDo+++rpdv+g7/iwsuYKZy/WiDD/N5V3wI38vjN/vHBVR1JLR
j+kWekHAqap/tuHePAxvToPb850sguHUtblSMFKOnCbcmbTjG1Ugo+KK4mDQb+v6CgbhCSHXQkU7
CkTPYv0Dca3y/X3aKBx7+PQFOP1uPUWMiCQjFTsF/AmpbnzGAA0F2jorqY8Fuu1GnHKlH2Q+7sB1
TBPDX6llrzKcR7fTlDf17ASMIAxz82BZhe3ygq15Ez10HdPFlSgH7a9CxPgMXQET7BhnKtaboRJ6
oTcCt+uDlB49dK4obTvL/SOCMX2OZXjP3dv+TLPUuyy35DiDj32VZv1ZoHAJDuq190wTihgV3uDv
iNjSzPguoJjevTncTnXwBZOpKpD8y/i/ZNUD8/0u0F2QtMDWLk+yODQZ55Ud2Sznd+jNZ9zCaoDY
Stnzy/SnlYayPDGOcVNU6AnbC3yGG4vT2Y+/1tmaV26hoo5OkDRTwaz/G3VVNJslQNWl3otgbdU9
9kz4RFzquE+8IQ7fQVn3YIglNoUpt8YWYRNTxPAOH3HvQ3rULWMQksVRD4UfDlOA2JYVP5PQCT5g
uKU4vUCdV34tOo54gUs/+eDTqfzrtSmfgaAV3uztf4vKGy0hRjQeG87Nlj+MEdQrq9FBSlGIDOPn
96kpm2/r34xSWzI00bL/Ah2gXTMrN9fFbNzTO+dLVT2M975jcdDCebZryAzE7+vlthcJIdNc1RbL
QMuHfjou4DMwKDjYzTC4/JtGAuurN8kwb9TmWs55DAZvBZXYxPvoAqpzMoZugCGc3r985OX0YBEi
5Y2XXsGwayDuH2ssc4cpqmxGpvBKnV2NxDPahazsflP1zVquyXHrgvznf3/Ctan7sbzAC66rIiC2
5i9rgmZGiFhVxFIfgsku6H2PmxdF9P99Yx1kVDY5QevZcR3EzTaepQq1hE10NI6zZ03fUnmBn0do
xKcMRZ//hva+li30mPAT966Vr1lKy84tPLLlor6618X5CqmfdxCZIOI5T5yA7I/tjjEBVpp7Cioa
Ge6QuehYE/l+ZSepQj4MKO32SNY79jFdn1BS4Tu97Z96ImUlWlqzRwC9xdtKwXA8e+Fg43xMuT5g
mDSPkWbl5atESR3Oc0gUdYzewnkRQhz/vY9pCUdIezQWSUinhEH5/2bf5xSCsm+79Vs1KusSJWvx
pNyEkEmObNdaDs2qzUP98Xy2Lac2YVK2169RjWzT1uRoO+car3InoXItSstYv95EN0aUUnwKbEBf
/ygwStChOjWOgksw+eMVodaNCrFJd7VwqIUcNRh898Gl2xD7HM5L3DVJPCyA17tZYyOnK9RlKwSq
IvuX/sepzTVznRVTvtZg6hSRHIfYv0DXOsXjjwDsAXDW7v8IxpshNiFwXyC0SNZzN9Im75HhT7Oy
BWXFYFqGklP0GclzbaVHiDJdviKACZOeyuqpSWGYFJM48czDuSXZV3oyoc5JK/80BnXImMX5lDr6
Gu0tBKByPgbNFlvBknFAaWY6iuuHqCCBEafMalln2S9QF+nkR7xCGSdkLywd/ZUdMCq7l4ocL+/9
3jZfANMOSOPdV02+Ruo4UV3q+X7OJWnAB5KWcE7jjSA4a6MEyyqrODksvhM2qPCmLhaymVktDnGn
fgHtCa4J/R/WgEOpg2tkSXtYWen6YaFUVVxA6Ioltjl80WZLus69ZU99iJQcLDl8djWUSHpAip+0
kYz9dTapkjUYftYSRQlLmQAZhfaI4cGPPfUv0BkSL2t4aLLNZf0rm1Z3hMpB0UEyXMm707Nc9rGm
Dxv+0dEnLPT4ZpjPPODz+9MJdRzFwgp1T3vQp05BFIpUFbuLa/0ZJNBSK3g10W7+zXdvqTAstQL5
vJ9nQs13HXLKkKQjdyK723xLn94Rd4f4TmDSZTJ8pGVEtkxnsnK3ISk5HUrl5L7Vy3W8DtldA2Y1
ct/trTeQbbfYd4evE3U9lGLvD9AeHC4SEkhOaELgK4aQnoyyT5YjOsYvtCuHqJOXdX0Pf+GPdpF4
xbjSmmXfclNvdaVWs/iYZVJKasYGJTt06CcvbpjVxVNK2YnSpqHzx1SlF1PhkzYzxHQwZR/AufNK
W3QucvqIeff74GP2zS01wqxzdeExxklzMUNeKhu2N6RFXC0mu2q/0j1nntyd5OrxbjnHKmxYr8j7
sV99RiUuRKPFOccVDxQ6y8Q8WdgGjP3XaINJsx67M7/wzLWuMCgIOG9EYG0psM8PiI2/shv9KO9E
ejBTOq2JUj4NrIJnVmyEHa8TnJOLOUpX/jKI3bKuTbu7+ft6hLEw8+dfDhQInfRbUVbmyKDSk9EI
QIzcrVcs7xKerPdOq1wPi53elWrWUD7HCt+EZOFJDG7dbvP+HobzpOsKP40BTYcPHwcJ7SC7Y9i2
K8NZz4Uj/0JUn+kBzI7zoL1JOzRIPIu5Qk+M/Jm+UdDN2Z7bVP820yN8Hm099ojL0XsLqowSFoC1
8L07WRUWTHZxqlGLWFUXyyr5zedEF3annu7EhDsuuu6xMD8uAG1q7v2zM4SQADf9K+KCYXBsTj4a
ALHP0jqdIe+Acg7ZxQVGF+Dasid90Tp4lzQjBAzXtV88I1zMaLH1p2v/n8ItGAfmXaIKdATWymlz
CvZPl0pF9lpDBIfA2KhjAdZFMKP7fUUz+ja9uL2bFGrdwKo62MDLh1wCywXEkTkrffyW85zV52Ho
cmZLs4egBok9+S3Uxsn6iGuo5+9YJZGXH5rwKtLTaHknsurpIhY9d37WFjfmQcZeBLUQwXy71RHv
UzxT9lVJ2p6lodP5g2a2e3VYtw244ksMNmwst9/RdVusaJoLpd5+/5uSNzaTwi/v9liQ8f7JqX2Q
ISq+QNWp6L4Xm6I3Mt21X/lBl4OWaUdehF+xyWVmFN2hoGtaNeKhUNWoEoxfiJ6lXKwp9zszt1Tp
U/FRPivJYoV1tVWwd8LW0R3tRODIRPG/Ux/vRS0q7e2NDHy3Xfs26X6Qf8ULp5w8JA3pVhH4w1pb
dO1dfNeeVqhqu2jlj6Rlc97Ptne18kiG9yTGjhlYy3SnrX2X/U/fTwSgC/dNCoZrWigBOjHg4nVa
gKbIaVgoJ2njUHW9im86ojeD43E11OwDMpvYlIILDtALTB76CW92eX+2qgZxyLqf8cI8R8PPA7MP
HRgNIx40sgmJOLJbTAzuILeaVfkBiFDdzqo/QQI8CB5fgwNLyBVG6G0KxKdnh3tOcRTxl9SkxKbV
WTfeu8L9uInnmLuI/AMDxeEKSP6j3cIT71Lpae/+NLgausTa0ackpxXfSBd94hcsRycQys/kdSAO
u78WrxkhykPP5OV/G5vYLTDah+ReudQ1yVZe2L1+Ask0kJ12KHUhb4I+mNUsSGLji82n6cm90Lmm
HwUWotU+ehsA5j7e1CAc3DH1CGPpfIJdyJEXriMx4QorVO1w6G8d1VUuUVrOUJeW1mq6Cqabo17T
37Ey61eRGqJrn+0tzwZuZJMVKXQoetk+lsGML/GK/RKLGgX1KdO+4FrALmC0Rh5RcxJ4lH2iHk6g
aBeo0sWbGHWCp4K3fV2B374YN7hesppfdweqLRcMmh2czYEKH/iDS+lYOgaRGQEQeKGAOYQ5KIeJ
VzCY7d1HrkMddtVLLqojG2zCRJM/0I/D3QVxpexr4b34SUiM8r7d2gwcqzQbkqnGK9+mrXo8Vfiz
TpkdJcH/zlj8JEtdVUnsljvrSpWZ/C3atHhGyu6aeLFjXNKn3ZgFzF/metMyaqVoHxfUx6rJA1zV
hhcgVInKHQIeByfTzkvfdpD1R54Cp7IsO/xYLTd3l3VxdOkr7hIHunedW88D87ROiGUl7nnTsl69
lKnDmgFkIuLG7on3B0qCk949tE6SF5rfVH+VDIkV2T/LWKms77Pi/XN0fXs1LUAlIwwFyW3r/W01
acMspsO3noCP9sKyYikrXiR4v91mpLcT8arD/PtH98iz9D2igt1lpjAWnzVXDrhIctUBKc/hEGve
znJRIXWH8JucfEmsqKyxCfJwFZeZHUVMHw7CvWJegKWY6ctRXb2dPxWxMe/qiB0LEFIglumayyO3
IskC/kYnrG4yzEZ57P4fQdT5ZIm662iuRIXypWsa2XxBUhN3Rqj3E99yXIvP3uxK8IZKOyetC/LJ
zLqIyy/nsqW9Yz9h8cZVwgV5yEWIhn4HFxFtstVVWsuIozxacbal+S4YZSxtIdcLDVgCBAGqXyUv
xoPH456kB9Ojc0aevli5Mk5hnNCtCDUXbCSvsY0xm/TbGWZVmcNXmOE/di9NQsbW//K7HEDYziT/
gSaVp+i3j8Qg8oWUq6oh4kUGKpPM7Vzhx64tZ0zx6G+OMGsSerGzjL1VT2re6RMi0JZmEub1Xtyv
hHnyPhb4hLBVCpK15ZePWk47XfKqvE2QsImL8dSSX7i3qVUjsXn0N9vjDqLx/tIIEejeTKxd9Am4
TVh7dyDmm9aFCLInTXGYko8Ur3Rh1TnlSdF/9ZuoyhBNHyrdskToPfNF2HNILbgwgXz4tfenQFG4
L+WWfj15UvD3t74tFuNHEIr1bbIgI5HMOnMXEsTvwtIkO3qZvvDhDGtSREBosHWyeGqjEWcJuVtY
yoxvDfWb6FZyRjLh0S7sSBXCYmyhNfwX9J/pJrjuDC0YlDuJCMhMrzVUlrKaxdidVt5elAcP7zfL
gu/GEDoQMLttJ/QXmqE58khBqeAksB8lZF8JNDtk/JYszZUhgKjuKSUuCMIQnP1GhujzXPZCmx84
qAmwu6ClHd7Tgbb69RhL4tzHzxAgqANMNB8auuT+IVAZ2zgmvaIGwWnf4tRAgjgejZTzJVRwOlSu
bWyKVpMiWxpP1yqFZNiy6BN1hNNpQr/7aWP/dh93NkKqtItdaLBuZ75sq3nRhgUZntlrLSYieLuk
XbPcKScNFwHxXmoJ75vX8IUkfhsh0lSe9BZdGRoKV/TUeHD0Xy/Ww9mkVPSIEtLSNexHN8TkCrOh
7VmqQky8LkJvqzwDcMOBE0QmjrXCPq3dYExoChz7KUjfNQXLy84yDlo9feJphPhtC25af6r2VC5a
HYKr90kzzGVnEGpOFahSRHntdZuQ4kS/SZvv72JEhO1SD29m8LlppIcutJ/FBqv8Z9BWFRHt8dsk
csnaler5mYgqZOh2WXK18NsKt9D1t2i8iuotPeWVPuHLeJCxc5l2M+16SMKUl3TWzWa5yCJ947mM
Q3kLFl1CYn+lMWlboBNxoGMC3+inM2yoxGCvyTfVhwPPrUH3QblGEv8K5H37qTL2RBh7IQQK3JVG
Duz69MQMYX0vQSTU/GOlS4rDxTjHQTIz/8QEVk9KEdQqyjxByM0SC3EiJCdUu+vYwDtXkQFGxZmH
0pK1bWAYGJJhPBDi763AwoqWJkDuFFdU+9jbp9GH8eH+mudE66EeIMXtSsV8z4SXAJO9FhDsGpx+
IS/avhX6CAIBBytSlFBAOifB2jIO6qtuGQQre56qyzOzykqlmiH3BOLLeAPcBqQIfV3WvCGqhVsP
dtiJcxXXtQVzAwz9Meagt4/on8LzlP9QSQgTMndhb7L3bTfGtUvvcWME4V6T9/espkdyCIU7ODrD
CMqjEt5rGKytUZredRAkLVWV2Wg1pc27QN5a0avtQc4LSRosOJLB5vqXatHvHnt+T/g+WyiGvtam
ctb6wljHlailHHUaIIZxIMSTj5Yby0BMGT98WEXqJmx4fw13LUv6E4899Ww5jMUW9TzS3bhIGwzQ
a5DsF3nPMjy82o4sYEPyv8qrAjtFErnRhFMi0BrmiUknQmGZmYQdNJMhZZlJ3NUssoIEnrDypoYL
DVcy35tU5rLQUZgIzWp9/5QLMPK9wwz7zOae9X7TfHiVeuA1adhYxcdv7YN1LWPw+CW8EPPw6vVE
SQM4+0DEKuT8cUkrhaRd1MkAs/jbUBAklj6UOd3UlqxV5IDbvLfDVlBuMDH4BbjtXbv2BC7uqrjT
AXFMijspD9Lik8nkr8uFRdz8Tzd8KmZW+976hGhbykgjJLf4Hxz1dl1VWtUaxdBrTe3Ftoq7nsOs
9gz2CRBNTW48V14XclETBJ5KFNxBQ3VfWr47694YI+GrrwfliQte1yw6LSg4e+u06Yhh2YVfo7pp
FFntF9FMRhb3O+4CrBVEPDAHMhUgrEPWXZAuC192/+B0tFl0Y4dgxJgwKjgVwbIw/k04RKBOsEDE
LxZmT7gQM2OoAEkZoGiGvj9ne6Dw6AXX8JIlFWyFfT6GqLBMwdWTjGlZZ0T3kDCniAyJ70g+cg8S
urdXTYzZfZpe9j3aIp1gf60gHeUlI6Me2BKfq+xdtNW6KH7iy3/+64qJp6QsvZ0q31aEJL+g+AOH
UHGTFW225HpetpaMhRvktdWHFMJXuxx8ObTPgXDtuuaDebDeTcbEYQXjiFOCfalmsbj4FmHM0blO
9v2vY3bol/n3xZZs06glEbIX3Q8ZvCZJeg4OYr+ou8XWT2ord80reEl+YqcSRMHApQk0GwaPeJ12
fSF2H5nevb6BNhaB+YR+xi4zwtItmnMohl7c4bm/g5SasjSuSpkoyUAIcPSfbHoDcym3tBWiLEqH
MqWNj/px5do8IXrdb+W5n5umrGZf0VvMM36WtxAoeSKpgjauSovH47c6I/XcNqSovtzc7fY8wsiV
k42Y440VnJnV2RllOKRpCp44lrxUDTzfdNwr6mmGZkYX0BYtY6d4UiDkBHp/QotWt2DnfySDG0qk
NSqsNH8+///RcLNqolepRoogU1N3eu0RU7k65nMcQRCkmyeHRPsshta98FJSRmO/W9Bu2a+/swwB
i61J1I/DZM1IdtDWdcqYMP5pFGvyUDTAJb/3sbUFtv+V4zgHN05RC9mLMYJul7jsum/A2WNJTiMX
x/CHQah7Ona4Bigg/5luUWKA6u7UAFxUvot57f0USi4njlA6SkvEKkfccc6VUItv4CFFeGjwVmWd
sVrymo9igsL9EuMSTZXQGwgaO4J5QvZHbaHLKFbNQqc1wcppxnoohFRidlrQL/rCQAzwfbbOwWs4
Hjinpm0U+JcCbBXI0Rgse48jLrpmthQyaiGanLS090fSCDyNVpZR/wxqNcvxUxMepk4RrZT3oadx
pSLVCj2e+nswtm3QVOwn1DATJ9f7GIT/B4U9e798n3NOCSwIwLwVNtlcZeqT0cRb9YSeSuehNeJg
D3upLq3xXcWgmxyEqmSRm+0Y+SGro5r6OHYRSBPL0Us9baZVvYGC30cpFMRVvW7vYsWfQVtq1Z4d
ISTNx6FCp/JZSUCR43IpWx/tG8uZGChGho3tBqa9Cp8T6q9A/ZGYnfzx6AWEP+Qjj81XcGJPv7A0
NlNnH5GkXAr1kkeHmboR/GJaZ0VaB9gx5dtbglGZdfPOD7LqhKRkOACZZwYsecMGSVMZRLICIY9W
rRVwQn+VZ6lXtBUAr6wWR1M7s4FCIiYEhjgMWp89Mwqpc+trgcmzrO+Y8knq8kq+yqlsZd4K/wBc
srFkOFncqE1HoMfLSYJ9aKRezowxTeD9OPnMwr3+Jg5oluKKkLTJ9mWG1+p/vZxIi6xgbWFXtLdl
QuWDLACTQ6eRWq1FGZAawLMqDtk0S6mU3BOo4Y99GGNeVYn2S4Yu9a1h6nR3SoGbb3mbqFPlB4j4
p+EE5dgVrFz3EXvOa7KWZRC0IFRjahH41JQhEISVNIQHP9ioUhClUpInFHfsyqZsFJnHwx8k7YbK
MoML2Zg4ojl70fZpVSxbzaWT/Gete4yh6kto1Dsv4k84GjAyr2sH2y98G040AlPDnHqWIpizz95x
5zZI4JxMgQ0dMWfQnb9jxJNbzYWDCfxSR9mWNDuFO0nWP1s8jjQfhdj9bfF7Pq3QoDsNz/8mgJzT
X7E2hntlTKP49ffg4mxT47aBizqIKxROPpm7oK78dkJ3FMItbUnh+6/DP8dvO6nPcICQdsM/rxVL
0Vv3I+7ZtJ4AxT6gYnZiat9VtUvT445F9Ye9SwaQugQgfDn420hkl9EQbw77bT0CDxO9JE3Qxweh
hQSy4duiBfHeF7T1ZzKZSaN7trdpEx1DZeQkgalsUPwssyCEAvFM02fihNspMyIYosQFsg4I1WIX
BOwRzC4uTyz5TaqevM/YLcjSNV4gGhUNy0prANQKJXfd84DzN234IpjCFdrTntdE6mwJD9NVKZAh
abEldYkPotf8oVMpqqp55D5rIhyf0dX+VQMZyxYkPuUBHmNHpKpHAJnR4mcx2IdGvasLUoftuDAt
SFk3RVpeemWMaitP9tSO+TZVoMQbbBYVgFKTgE5sLCl7pxEGwjRwIEd6p3Uudqae85zIpwG41/mB
bL4zT1rIyFXijIwUTn/YmA7zFbWW+IXWjQaq1hXAsThfaLv4MmWbrFTF0Fn3GRSVdyDPSki0tKKh
7zq69kni3AJ/caqFzwHpHwMlrgHSggiC069FsrPs95RgGHbSfhbE2ZCKVW+fTGTObPw69ZJ3Ia8O
8NorN8lSaBWm5Ze5byHHdmK1dGAF/sZ7C3ewET0//HYAtc3K0zj1KLGx1YbP+lAhEbi3CvPP8JkW
gELQ+iz2lulDJ1v73YmIcTEZOBCWgluMB5I3wm9TaQUlMfJ2VrUshgykRRiG0yB2HHd5FeP39ZpV
bY6cJtDcrUuNsW9kGUEZ+QQDBfiGKISL5D7ogK9/cajwDsdkH6rLJHavjhMvjmVmVoodzA7oqn4G
akT2KK/T9wciWWCwSiwHjPlXJELIPiVaV2VZr1Q6TpogpaWCbJDITGZkrkVpAToIyVBb3tafnzEp
vUa98MOeayuBPYYi/BkUrcbw+Q/98beMowyVsWhJBETpKxWGhzf3bbIUErlnoxTWesQha0ETanxQ
s+f9QaAamIRn0Tg1enmJzKI8ug8uJw2UHl4oi55NLiMbZ02CWkbjx5WOrNMEsJZS3cbd2vIodzpp
IMfaxCQ5FYzLIIQG3VKIrhT4TfVipTcbJOxlJbZw9gVU1sONTT5sCAT+Nf3XMKuoz3Wxe2TV32RD
HIz95YYZgMLVOPPtY/jnJiJGKhR+dDhq8pU8Ivw6f5AH9gtchl5P8f380SjSgXP4ikuY/N5CLeZi
9cGn/RPoHQkhNABOYH7U2kZZf19fxxYGqHNcZl1UrqBd5pAz98Sb56KLRP3avfa8yEyb6b8UYNFH
KDfSu9UMgr5dDfcN9zU+1Ma1iwSvFDCIZbyJq4PrmvHDSXGmtaA8oFY9Cg0DLfuC5PRJvFHXrjIH
aEbsKi/u2E7n1bhphGNtKW+MCldoAYuUrWUsXfP6bmeMXYIFNjeGY/WRUcHfbmmi1zLRdTJC13wx
/8sefKf6mLvNt4Y4c9LbR/z86SbYkFV9utobFZU+eygNo1qqmIrDu2omYOJhIuFKuasEoUApnaqJ
1EHI9ed7b+y4OVpfeWFQu/vE7Sc+jVEa9LkAFz8ySNs1+h0Yb5WKCmZnKJvQSw5RmCZ8496UloQD
TxCAtN3rg+Sx//Iq6INehZhBbq7QybqdSkHEAGH6x9XRsU9ijjZLPWaQtfIccJHcWjC0+iM1Dsym
Zd/8qbQowLZtg4MrQV7SgE3puS0HFaTN/JUQzAl0aC+7j5guxdl53UXaZFz0RL9gFM0Vx7TgSpGa
vV6o6CUy9fTPTz0dayyRdywX6kUSTC3loeXxGuyK6ru8ZXa5+73G7R6IU3aCVH5OuAey3PmICcVg
sx4cqFi/wnqgRKrBQKL/HOB0fpt+FJOW6+9lGH2EMl7oOzoiPCmtLhFMrT1GuRm4wZVYXkwg1wAv
1svc8GsA3EEYHf0bu7jgp3S5Jqi+W8T7+2reFY3hhdDWJnrFYJFEHa8iN0+xd6w5WZPGZLT/d+3k
Xm6/nTK4rKHwyoHFAcGevS0CGDER4FwiFtm5VfmQHj84fnmxNsgX2Rn41nVITS4TNswXcUryeg2J
/qXaEZvo6FF2X2kMVHueX9ZrybSotnPanz1YPlNX1jSnYLiNrhyn4DHYjNW6Ny4OHm4pJ7Qdz8of
L51Cu47xawg0wedHiznsLidBh5MEdr5O0DTJ4+A0rYrwrr9BtkP/5mBfe/HO8KWF+eqcBuDGIGd6
Qf/C82YJc0cUIMw8PKHtN4t1DQV3A5D0eW34nnkckRmV0mqw5jPgIJi4Z+OdYhXkk5Ou+O+0OX+f
Ws5W0r3b5XfDUsMkpdekdJJaTr47Q9Xip2VvP+DIGfu92OnnUy1DCkfjdFPbY826x33/M9ctuNO/
7TZAif02CvZezQfAduSJoLdJEgHJKMsrHvtfFctsoxDh0n8qG3idKlqyqEi/Az7TOKiorXIflIi5
SZGSHbrsPbeFDCtKzNSadACIx5rYtdqtAD42gWRpw4+OQpUEJFLHUtXA/JUMQ1K23kBVTtYPx8xG
l2Hch/Wg0Di7ac7qWDJ7kE2Iq6ZIfaXMoR8YbdViRo83gnZJNogseYf6hTEmR8Xzgse4eG1y1jkP
GBT5v2kSumDTKP3fKtFglSLwanZHyY8A9BzKw4+gK/rsVo35ireiKVCPuRmoMHDm6yJcreFresSE
YHPKCXFLmv+oNchTfn3nOf/D5yA0RNtCcIUuWzJq+WBFqXGyKbQ1heQJlHy9dkzbDyj1HxjPCaXZ
ApPiLOTZ3Y5fh/EpQhb2x1cPrUTb7PdicSxFi9rnlY8ICW2l7PlkWumPGedcR0PAYnvbPwS9Tm1/
BXyTwzx0alWfLD6Sb+GcioMeyykna+VKt/wtbB/bfP46oBEbefpbcEQE58WLuKGMJ/VMqB71jo/j
rONZvNpd7GNBVl9nM1pW/dHWCaAdtvEP4QpJTSlCr638ea5ylUl/Ms1AW3a/XyFSdi+AZUlbRIpm
THoFc8zIjrFq5aLUECdj7tbai6OYhYcRVm65SY+o/5BDqaxGGXeSS2HazUA77Ao0DZmgkE8fxHNp
YKl8n/aVWbZlrImsQTZ3SCTYdILBwsIkNVeoEnBNtf6osUKFleAtgDmiYdYTCpXq9D4Kwrvyy6TS
vbq8rNuoS18YBcc5CuCUuwJi/jleusUx3mYQxh7sjWOS3uNFjxNyJgM224VJg9sNyY++a+5JOZbj
Ea+Rq/r5R4O8erU5su33ZhtsRUTlwgrnhwguvfd0H1wedggkMb1rpFcqUKnEtzC5n0UIQ4D7TDVC
7eJ9eAtIL+296/hIhKJUiehYCrGpPGCp2jOip4t8ApiMEkrRLk6oLuglzYuMITzMVHF1N1bCvW49
o3pbcy49GgtMVmFiXQim9OwLkWmt69BU06Kt8m9RI7lX4kEWVeErC0cnMNWYZF91oS6EM6BJ9pgj
kzPRK5Ab3e7Dl/U+QOa4kl18egZR/Ax8gM24PysU+Ev5IF0gKVyVf48X/fwjSqbYrqWd6G+3YNNz
nZDadA+e3y9a9O5XaGNgrGykIS5UHsegaMRMSul0whhyvfHYmLubOsB27jOZoDWuVGaF7WbEyBVq
z2F3Vm13JYwrFbGwCj5pdHmF0DZcZwaDNhas1lbqg7b1o51MgrwJA/KJorwVUbmYaCEpTtAbFcsT
dklU1pT45InHCe0S4eGc/hFiCj+dalVzE80bbeqdxSjx3ar7Qg0V8Ch5b6Eo0bOukH3D90AQjx8a
C+4fjHLGxBErFhI3HuXhxxqrwU5sA93j8cuBp++zZGzAkqvlaSZlkLwEjKVVOJP85Rcc+4RpV39o
SK0986OFt3wQZE5ybjkQDD8H1LPXQI+dTV/DBGavJwkTbWNGNVVf3ghglxRo6iVSS3XMMTIZ0fc0
2ATQQeRQAf62JajuomuT/nsHlspaP77oAjW99xszMamWD58SFmkkVDj70KLXLZn5dA38Wzhfvamm
GZZM6EHMUTnxO7YxNCUq+CQ9NOP9mRgojFcfE3NUsdXI69s7cPOSCkEv08W5AwqMFVwoZ0wU+vFi
uss0C2Aa+IgjmMfMNLfd8ZORINo1yu+14ekNyXESuWUDK/Qd59UdmS7Tkoso8ZTtKQIN9B6ClvJ8
wmAysfzsKpYIChmPzkQeTqVC7VzqY6abPUOjq4lrTmg401gbb7OHCEMb74vcT7n3dVlE+/RIWezE
x3bZ91+uQDL6zXzM2TrH/ZoIMLjP59SRL6KkAfDho5SIMK+tz1jhltxlt08GomVypokeBgCRovtW
O6XbP1jI7j+ImDIlFUNy1nCm8KoncvE0SHCqNC6P6V5nxTex+jCGRkDofU6xnEueGDVa0Jt8lKzA
y9Kkv+4HQBQEvOcL6U8uUZNCyimWZZ/M6Nrd85OdeV33nehBPG2LZLobv8HKhlJUG6YuQoQKbvxE
nwAIBmgapztHtH99kkCKtYf/f2Lz4u303hakEbG6E+3N1cHTizJMTkxVBzfJ2ME3/+/SJZIZBY+v
9VeFSiOXTSbhysmkfyX2uTlFS3RX2WBamgSt2r8cYcBsMmR/U3tW4q23hPmbYcUw7woj6Wts4EPR
li9fDLx0nZMGVAxcLgdMvW6zA9yesgIhyN+5EvuzCr7Ka2k5J5N5CzSNho/tCEPbgNHoaEH/XjSL
saGhK+yQK2z91mHPclraRcECY/lOFz82M3x5U/EYWv+P+AbbiAEclfx9Ubjjfyk7L+oMpEznKfko
ejQ2ONGXMVE/HySirayxJKfgDPW5gFDFAoUZxduN/OFMd+RipN+3neDa80iQvkOKoIMZNFyuB87p
/CmP3D8GsLMlNyz3uBwxixjkGuHNHN0ICdHaku0u8F4/gS6Mhp/2Fsp0VawzxqcvxxEFDB6STSiq
LDtT2ht0OhVOERX7Cg7THeFPs2rjeqlW0eysIEfy+cTpKu2RPjqRbCUstkMZFpmog3UImRkGw7bc
wUlYUcrDpsOTxZN0T8ZNCP/vgq9qbdVKSFcHV245ia+GKceWq0EwvqbaxLIvzIhEImKRrjWkiSVi
9Mqk+AMempS8v4zCPIJdZXKNmAO08SnYRRlm7aykT8YC6fzl7XEDpAguYQMLLoVdlcsvSZTDR5rX
0JbeCeYwPtJV5dSKj7x10GAFQNxI2FpHPJ1LG7+aWa1nHNevOKtaiGdl4w30Zc+ZffZcxTU4HICV
Qbsq2LOhvuWn8Wlw9guSinhYUIlTwH6aLEt5f69Sx7UHBGBcLJC968eL6UW2kCEi9cFpVNmwyZ8V
6WlzkcDtOJouCZ44GLm+nJ9ySrcus9uUjJ6likdSRasyFZt1ehJqX8Pp049zTI9nIE6PurzmBaVk
S/T+GDcpYLWcc4SJZupUcqmvDpcSEOlNRXS3wQLFk9To2c962Nq+ExOUZFpT5qmzT1YRGr2xrx3C
aEGVvyTCRWD4NtlBTtzTCj2Ak9qLYDYJ8hA690Z/ZPk+Bc9hUHbUHnudrGPCTYSsv+wQ9jSzQXuG
njxvteW0l6TXzwg1Et9+DwUtFujCxC6WjBooBY1YnepbmP4O0d4iHdI0zdTxonSEfLm2+pxbX92C
WPlDz9NbqFvc7M/xfo/eU8gvgVOJpnX7IvGHQVKxRXrtY5rFuRjXCyjyFccGmHUmiCXlIKgxRTA6
iGOljxddkj17zIpfMepRas/vkreVxc0Wws0oRitctjT3a1wCgeZi4OJr4RezrkCIBjgESVvPFcaL
VdMXP+F+c+Uh2z/Ub32LIOyDhMZ+Phe1PDXDKFePxANm7iX6tYz2mJzvfGcM0qWWxUI9J/MBRhyN
tpdQqub62YyaIlJw3OLID6ygrizvFg7TKOpt9CCWxwL0vBPCnVR/BfJA6WLJTppgzquDqo42D/SV
RTtfuzHNBGAIp5u4/1dHwbI/iMaCvxfiAF+PtLGfMnSTRjUnWhJDncqL/veoiWlcM99USXlmJBEF
S09S3CCn23JRpNrhx9/dPliZuWZEArWniA7SE3PA/66q8MEf5Z58tYRwv8UqrfCcoCfdLQR548Fl
EmEfbOJpKX05EUnBrxThm2eHJ2h69w111nz1GBgfgPpbrFsuYugjjSRbbg52jfVVh55M+2YZqLKe
RKKHZ0D46Clmy6O4Lo2m4Pd4l2AqOsI8cCrys02R5HyMJHfqRlWLtXRWUd5ReSx7LbyU8+BzGugp
fdne1M5/ie5Es5XKQy6dKhQAHsMYuQeYrjnEmZK1acmVv0wVCq1xJy5w0ffrs7m+eubXoODC9Aib
pqFwD/bEWff0Mu2SPkeNG33cP3shUJy+OVcjxt3MNU/9PwKPK8PwHU9kqQn5guhvawGHNHX9QPIu
Y7MgIC2ae4dMGqZ1etypbhEykj811CSQwqN4JKCP25mYks54pue3cJcuV8b0IIVdP11yObS4wWfd
2twCSXi6RFo2CfglB1igTuuwRNxvo/XCa8YM/nm6qz+R3V5yLzP1G2ScMC/mm47V/c+4nCbOObOr
9aiuB9BU0J0UnFpEVPtoGmCoZjeBkTRSea3D4fyX4nfxAPZVJsF2LjNkoDg5TFJc39ohlocw6RLp
naY81XRbBgWwBcZP7bUENyRC50TXP2+gRMBEk+B7RPOESxiQM2Y9gRgUkBZ0sOU2phUtF4hakjP0
hVBGBu/fEasZaPav/f8BSeQk3q4FB3iuyxZjiIM7aGwQ2KhCahnDOfgZE6jHsmhawxGOOZd6SKgr
V2QIVr67aowKrxWOAkyM7/f6CT0EWaYEFvFISxK1WNtkiCk1Cc6xG+C+zwWkyvBUDGEh2DDnIrnh
Sd04j4y3uHVP9GI7CTzXpzaOupqpMu7QFZwuc6DyH/eECkfHF3Nv/qFIfQS7YZjbZ0PE4tZHve80
Wmtu8GYaJfDQzvCHhELb9TlGY3mTYEeeIPnk6S0Sk+8pkcIkJ+48obbOtl/RosSkjlDrboHlntmF
8yw5xTrafJaMkERA3Ky52xZeXeQIeU2kNkXwSRNyogUf3C05PTAgWCtf10eXg+ZUJJRciZAuLEBe
TBj6NYS+RS41Lf0oI18LkzpS4dUrwrDE6cp4xMT8PbKNhbGZULV5eZToqAHm8ehufCcUANdpi/zj
QOXVIXhhEftFDscWNy7BxiB/c7i2nwk9thT38wupWtkutMi2JOpErEQMdp4yVLcE/gUm1JCoG+50
8JXPo/ceQwXpfFxorPc/+3Gt3wu82chG1sV+n9aw6BTNMm8e7WtTwSLDhi1w9oIuTDZRylxXT/xY
trXJ/Qjptg+50FrFhe5hCLOrUiKmOZEYNYSzXwkf41oIv2QPLK2XXNfya2ZMuyxAC3AHTn/9CCVv
SnEX7H19AkztXBBuy9v2xYv6+3SMUxmuaT/HwBUTUyGZPf+mbKoOSFnQ4e3B7GTztzz5fC+ClLnz
MWIorvvnovCpfLH/lj7jie5pzp8+yN466eazT8X8eYAfP1wSvgl4uBGyQgLPn+KM/7MeETGEuNgk
RYl03sRM+byhV70rSLrIhxTvztJizJwbmq1sYXV/LQ8mb8jPVBTtPqNSb3RDuU7v+2+WrCgrWPDx
HIRThouQY4G9oJJVn7RteEWLTyyII1KxL+pneMiaUoWGeOZpeiRwEq8BmCpoHWky7vT0agEj6XrG
BjtdmxrUBpO8a4Sp4iU+WBH7IpLxJ6Pa7akA0PHRvMWb3RMQvflto6euLwEctaTJ3vROHcK2Bd/s
kNcOnJoqkN15/C0D1BJepsdcVgxJqvFsl+DFj9rCrtIaiVpHKpPNAtOd/irq9WBD4KDIgfO0jJHV
BdDiz0F/yH+I8wYMxYTH9oCesWz7avGBXgCOFC5T4mwL63wA7qbw/h+tOOTn6htVHM7BkHl6V8K0
2lsW1USx1v5a8Dwl9rcfZFQtu8F7p5N6G2sfC4bs+aynPH8Da9FAriduRSXq0FQ37TkNCrz0wOLf
P62WKYlLqSkW2JCGi5gZYWQNHzPFD3Kw0AHw0NhRxYaAClo3z2coA/fW9NdfzrLymdVycb0J35dU
nc1ebIUcJgBogurH9MFbIf7ARs3YMt25WzWJVSIM6W6/TShWgbcVZPkLu/60qRsO1TWTlx8KNvt3
aN4wI3iEbNAGNGDsUxirfK5NN11YKLanIUdEXLlnezLBaSo+lh6MqFyyfyupwv62i08AWFHyDiNs
SOpq7zWM/FOpvKM+0w6x+hVfZuHRE8IOSd+5WwSzAMnFr4zMhyFeOGN7iY4fRB954b/ZEkGuCbxq
XzsGRQOFHR1J+TC8p3nKiBTMIw7LreGo8jAAModrICY7t4F4WtAdvWerHVcAy88iEATBTDr+G8Q2
8QZiEGVGr88lBMbcoBPpVIxie/cQe3ktwA2OytFwFJSjNpKjFYLnOfZWCyaQ3SHjEOsyTWlaPLGa
/INo1YW9aC2BJ6zKmRyEcx+Pmer1VTU1DJ1kY4o4Rb91ABFFIeusL4WVZqX/cnpTJihThUyht0TY
pPalgzfWd7RcAnek287LmhLKb4dQX7REap9DUofTO9XSbGKf98Bqtie0rdSR2yin1AB6vptibwZb
wTgZ9pi3WHgdoWPAVSfzmHZKACNLxukVWiaDZ6ddi82xdh0ICC2Ak/+gTs9cz5cbtehvies8dnzj
Py86lObldDna79zlGmrMfQE1szUdJo2jjwMQl76NTec3GMp6AJg3Ae8BDj9tzmiLGXKAmxPR5x3Z
r1wOUB0RMxaMjoyt5x47f01H8vUXDSrKycvQGmxE9b4XDBUQ01SLE6ESyZyqRsJRiRdjpw8QOay+
7BAIUece/N+DzIvJes1e/QDk2HntuED4YbCtPk5gW5HEVrczx4gQU/Hhp9UMffsJuv+TNGgQZRQC
Br28L/omAUc8G3tcsUgfmWh7ql/CfxB5wkHzuM+VPyoJs822kLdKVcT9/Zx0eIXDQk03mjQT/Ruf
IVX7M0a3PprUSzudK/lfwLTG6E0cH3VpiA7bOU87sQq6Hm8YDdoZb9IYNyO0HSLxdHkhC5qRi7nq
v4lJlXnEAEW7gyK+w5tbI6Q8uRiHpzy+YVuTCGz4yCS66f/mpE3k14m5XXKHZcWZX0gs57UAzJ+K
0FAQIX8fmWkllQyCBiPNe4Z9ibTAKtOysoNmIt6dAGVUelveKmOEEuRAMAoUDa7yWlMvDZ0J26JB
NJWs74ftm9tyhq0sCWqUZt2o+JsvthgjIBy6UOAEKDnK6qry5QHwBSTK7J/9kF96oTWlJEYgatk+
KerMVj2O4bXLd+m22NrzKoWuxxIp+2wsGbeL4EorNxPxAuELspCoLN/TlH61cd9rOBQFoRTKhPko
KXBsYWURwDQNW9oql+K2ijnyWRnbflm50w/se+dPapJcbVjHN9hEwewEB8jMjG+IxHL9nFcYFvD9
riaRF4gQq4p2AnAXMmdOJ6q1DrETnx02yMdYuByFl7e4Gp0B0kL2M1UFCtgzt1A8HRalxKmWZZZO
yN+wQTS747cRPrnCgK4ZMnWttvT1qAgoOoZjq/X+50xhWmxQqZii3D7muu23NI0ptmex6yz6oG/K
ow2Hjd/gBczQkrYqR9ffMVYyqI3KILj5O4WvT1901EVl7OS9CfwM2nIKpaMHNfy9pbPqUk3yMsNQ
H9+18iY+eTIPNlTvoGMbJdY2DmlzlV1gCS4OKi6H1+m5wRqKhM9aaUG6/33Dp5M0bi2txVwrX0x+
VV7ATh51Nu1gd2DNBF7/5FT20rbzDD4N2WLf14x/oj9RF5k9PzcDpgtr2Q+aTzZKVpEFqZdOB8sl
57/GdZYLW5fIl3X4J9340sKktK4y6h9rVGKy2I72xiAjf4Bszk5X7+dehyIZ8kbA1gIT8UvVwjP0
1qBvKEc5+xYyNVzTLw0clO3uO86RGwKknUx5yfENuDtV3aUNf7YwvXVnbRzKRVnPE6vVu62p9Jrc
8ZdJqed1fepc0wMdtUOJvD71hKw7K8SGBLEBh661nood2MbsL7Ac7NBB2VSP+W5IRHVHkARSPJZn
ta7okKWg93tSCN8Xwbn3Bnc7SPNLr/YuUUKBUAMSuXLc7mE+mkXWoSByWwvInjEvyLTA1onwX7Pq
eXD9JDblxK9G49J3afJ5Itje1TBpLaDrESG+TwkP2seNDlblFEVwNiM2lDQZM19X6UfUVFDj1107
WNDFQIrC0IACn5jdeOLLUbdRd2FYXuXLe+XC5CRYL6jIzMReLFh7yl2ydf4yqXDybtGzVSQJMYQs
dJ4cQWLYsP2YVP0C5nCLUl3vdaEehtcbfP/mD1EX5IDQq1Etb5s3ayKp6zz58eW3HvR0f0jLK07K
UeC2NGEDktTinFB7k12eAUnR9D/GF6Vkvn4XE+oYlF1sqQNWkVnv06O0zNuLt4bHUPqSZkaAQUpv
Jkh/muS1Y81qCj/+EcQeYLG2BvCvUx3DtkzPJ+lQvVLct2XI1C2dK83BafLv+rA4BXyvoIK6JddV
NV76BGbIWxCtLkaTglrWcoElKWmECinxAydngP7Ci7JYSWhD8YHKq/cYh44FY2eBtYO0cRdiYMpQ
c4YyX0Gzb86ij/bNri/g/ok2slE35jKihxADyaNa/sve+zdf4Go37A5kB9902FoAfenjyVof/Joc
oay4jPRq9ol6iGxtggtxlzHuNmnA8dF0W1Mue8ivkc7Axgdw5U6tI9o7VxiTf3VCP8Uu2xRgk+ze
s4EisPXS/4Np72YdiZ+ru+pBG0FNDjbAvnXvtoSv1RirMcD/UHrTEfVhgfdKd930nIXq3V04fvNb
gtc4ciq+EodI7eeTg5s46rDTFnKJEJOCt58K77yEhMARQGItfXJ0/xguIgrVT5xYd2lcvalW0ew7
GSGMiGK7vYuNJZFMZa19QMnkG5vIfBI8mHhUZAj+feGLx+9/NqPvyG78FoSI4t6OdwKjf+bCV+Mh
6a5VL2q5gWoEwqmZycxBI6p6o8zPg6+tguwNCtYFMUHDkjx4nl+A9+Xha8/IcOFqa/6Y86sUVoQU
ig8CZvFSanwyQuuku7pIiZSykyzBMKgzc9Ouy057ahdxsAGmUifD9d6lweXmBO7mOAo0mOkdyrvC
1BR1cX2vkcc1SNgNO5DYgfe27njwXc4YW54JxlMED05QevlN5KZ3HyCFB4ZaoRzZJjGVt1gdH0YG
Q18I6xbMeaUkuRTcEcjppCGl90Nh1U3etCEgJDURACAff4Zn4irR+/zWrkVvytnMQ5VhIDk2EoqA
rTaFWwQPtx+NNs/UN6o+aWH1ojvOt7eVYwHsgUgCF7gXGTwMnINbDaZ79FFAVksFYjXq5cV2nnS/
xhlaqqUzwAfrooMmRR5ecm2/G5vc9dvoZiGmKVLJmWAFaHG1SNmbJhzkQyh6heQWVfTkbHkn4/Fs
F28L4Br9Kvb+S97I9sqZvoYCfzmp5UgHVZ1ZKHyYAEyJkSen4UFCEEL8wmYKn9VwELqIzTrRZt9v
50aYlPbjU1cSefykOU854QTQihlo0Tg+jdTrsA/20qXcNJIBra5rNKDxwTh8kqo90cV6/I1cNDNW
m+tpK7JmqTd/IOBsozn70e6rNFfqOu2MDI1VXKs5cgMRYAoZnYFfHBhEXOtB2gQqcD+oklmIA6+q
CKnvpB+kCxTjAQwdpZxuQ++VGDgRoCeNMo9+QlANrdZFQBecWlNpB4WvdjA+l8BUVbW4v2rrJxio
JCKpg/NwPUOQPJZVms6j9szUurtUiGeVcx8lGHpvgNV+O6YJ1F09ki3qnWGvfyBO3TNnrkAX+aWO
yGk3BhRuGz0stQNw6VhdtdhoicZq6/NV575CCR9gIgVHOiAzszs64MY8dmqhYLzhUuW2keaUhw9V
+PTXQUrICop9Picpcj3iM3HXLYEaFrawt+XClLgnrZerIfBeG0owMZVl/pUfGvHiwtsPQHChGjYy
jBV60n7mgnXHHCdDo+4gtNtuXu7FhIsmf/cGbgVyJZCbkr8Na3SZqC4ym7mXxIdO/kJMqZjcu3Iq
ER85d9/CKvyUYX5r9qo7OwV9llvQKIME8Q7b5+ONAdxBJCkZkao34pb1lddp33YI8Kt+tT97ympL
IwlCTTfIrw8K7Upnv3DOnRR6ABDI7PdTNQXC+a0rOmuSrltYm5Sjo5QcHjsaykgUKEQop5qgTDRZ
mEoWAq9kblQHy7qRzq/BZjhA3TKYkbZKJPlgKgEL53EQrlQnBhoEX6Ji+izkNZ9ENWCYJ+7Zl3qm
QmW/p2mb+ZAJpYH1NaDJC56ddWoxLnoxPcRWO3h6NWuGcYOSA10Lbzfu0Z5yeKIIjUuN2xTg3G7M
/3gjqoyEpPPbgbjh6V83psoicmprOQbJQY0GJ7uuLwULyUg+ZgrR7OtvjStLWWk8gn6MzjJt/AOf
X/fvQ0xapBUhJbDQk1WRzL4K9nsdkLkTFjDez4wf7/AzQFjraWRVUrxlQjEfXP97TEpq8QN35i+7
X/g5C5oZZnvBZnIqsoV7p+04OC+Gdo5m8JhWNNdvFqjqmsSE1dixkp9vDd0lSiVhoArS9IQCH0YE
NanNrcPPOZRtcdVXCXJn7LzQLsR1UYEFIvUHMCCkhHmUyynWBFCI9cX68cLG+ExoqvH9XhKNG6aK
MvErxnnSOto/Tmaele2KboYF7pG/Qp8GRoovQvTIqyK0J7l8oYw9uJny7mv+LX/hE73nNm0ItRzM
9YpfZdebeysPp2MxwbN+IK1kDiMkZE6UwzFrdCvVKHDkMSzrhPGBaZu8p6UMvwh5mDvDTzuokW1X
7gxT4CAt//72zT+Z47vR5lTmxPnS+NTWpSI5/ZZTPU7ZtKgfqnRMBC7TnUGoasAbTnwb7LGnuKRu
binRIsJMrllzwKxi9ROIJwHvI+mZ3Y3Jm2GHdWyG+c+a+eFZ68sjjbjNxp0DIhc0k16BFKOQYTeN
YoKwJOGA6TepCn+PnS1rThAKWcDJpc5rLxyV8sO7tAbFoW0ID8BWwL1yQ/Lb+smqMgjWB5A3j09m
HzrwGM8qyClx+V8XlsparskU3b5ItYXHtWLyodi4vK92fl/FoF8EzrRK16aw1PjEOsM3cBfUcFQ8
L0BIOfW6pa0oHs1QD5/gOGz7574sNeub816H8Ly2Qt8rcgauOqhlE/dfJQESxmqgiqZ0An9qoHFQ
Rm+xrGOFyO++rcSOGxYqI6TchV60g1J0tLpYBskn5+ZjIOP0mOq2euoNYXR4MZ2DlYhnrzYgXFj+
QjdX1reV6D45/nt4NI1YI1HNq9M1ocG5fI4cn0eJRS3sn2GNB7nP0eMw3s7BlINL+aLvuUiRW2O5
QF6lFY/HdnsVT8Iz/bk+x3Brb/kx7j+G4qOqvDbGV+eWX+FkT47ONSBvVdKng4pUX4Ln8iGF0ABX
3nnzl71tjqEwMSrPDirinbIeK5d1TUSdT3SL6/N5NmbaZL5pMRFYJdxTgpKUs6j9yb4dZdj0GFBX
5H6t/EYmMRH00ZFEnt5BfZfB/RKaIVhuxqBrQsXS9lcrvKk12ZaJqCz8OHQfew95qSnRS5K9oj1l
Ni1wgPT3Ti/3M40bI7y4s4m59neg7VkSciuygzykks1nDs4F9fhHNkm1Gs9BgL/IihLe37AgnFsp
hhIpriNXfxNrfn/BHswlZHXiIbt4VhBaBwH6jRTWM+QHAMeQCXH4Z45EIgGDtObsqyxiftncHS/i
1KTjCcfeQFOhVFI2L1BjygE6ZXebERFRAKrUd3LSXkmOxI+S4mAUbBfH8e3TmsGYtzSOBJqeF68h
1Pd09Jn9lYAw583Yz0CTAK+f9O5dGoKjH57mFyqEWAcUKUaE9BDht/3vx64sCtC353iaYrXERBb5
ZF4Y36ouW1Hv+fO+QXLui84ZsbBrpTpP/VhWo2B0tasTEKWOfE5d4Bu1wPdfvxksFIkbCSNMV/nq
bAHXlPfVgfq5DjDl09vFJ/mpmARAjPkZnFtNA3cJOMktOjOau8dmwSRNmGCi0mtu5M5akz+96ga4
tV1l0iD1T9lf7nA72TLZ0fP99mDG56B+Qo4rcI6vyzb+R+ySarme+Fnzy3OXCtPdJt/KBdWGpCG4
w4WCqalHOkF79D2y06Z7CmIIU3Qatc9zCBFZV1pKLyv07qtF3TLiLCF5gdDlcPu9s87la3ROJnNw
ICBxbzycIidZzt7hzBd8Qp95Xvmyikkv/0nYzRQK3QPb0AWXnLQKQOA/En/wa2FRVxaI0TkvUuTF
TX2XQE3B0NtHw1rS7+qO2rKoFvqpMx73X0JMFuWrHbZP/fESdHmKB8yAqAxs9uYPdZxZa5h9GPuE
PAq6Dh/sC0GfiEVQNoHtpTBBSh2icTWtThe9+U8Q5pp2BaELidl7C8I0btPMqeWeZrkIngpUMNmf
WMx2LcQ0C4RKcpuaaOOfAU6mFUm7hxUc/XmVXg2Zsib8wPSMzDwP/9GtHTq6H+IAszO8w4Fqv7Ik
ZL/c6/qfgnK+UKBSr1/Si7Q8/W2h7676hIwP8noQfGsC0l9tqPkENti523vfC1i17XtrrduRc1NV
2PiL20O+xvAgpUZbzw37pDvuWW2RS3Jq7AiUoKXVnhENfo0kLeXTX/KcxtyXUXOi7R/Mxyo9Hcn8
Kf4Q1LmoTDPNBT+2a95x9A9cICI+gzl6gcxARXwAOaD9XhkMWdY+EYWsI1owF22iP2IRe2lbxjnl
07l/7QFSBDMofeuK4qjk6cfDxVueSfBr0Jn/WwgJsSXNS4msBmZ1RlXSnmWTxarAGngy8if3HgRq
Waq8QGczYZC/wfWckJGkBd/zubk8oVDBhEz8v2MI9TkurSM0vWlQvbF98JD2PWh5Cj/MIrBOefFx
XRp1sFfhGp7yHZn2zd7XMqnu9uJQJbGCMaHVnRkHXKjE5w3OXZWqxzQW1dpCEVu2MvNEoD9JOrk4
Z1jhRiT/S+9c95GwtQ+rR5IT4hofcfcqECtTrw6v56TlRMvKtlU5Hm6lSLZqHQkNe2+vbMj9tzpD
IOU6kIRZ1mbcsKBSjAxZkSOVpbj5uFmpx4nZyV3lOKZuZvyb3pFarbm1xJcHcjyuO7dHFRKlDiEv
p/hMJl+K4cRh9fRw4yoUL/yAOZJ8AmHZdhayIBZiBH1HpRf7UL4UZiAGIoNYLTzPa2uefsUI0Prp
mFi+d2Xd4r8ZSLdH4yMXVrqYcwHAHnuEg9MGUCxyBTmmkDEA21fA9SU1EKc9Pk6GobyktaeJmw3C
tURU/sZCrTy8urTRFFUOb3VqZ+9A8/hjm1OUsws1zHA6L7oy/daPC3hjRnKdR7A6L7+C6/Z0A/lL
Hyu8pYfIWIM+GcAK/y2wmoAoqK7mlH38zCLPVrord9jts8EpdviOYn7BWMy6xB1vXgkmvHQOVAJd
nPj9lqMhdpEdZltisfZKH5QDF2xX/PebQSysOTZ3mafvkAfhNhooj42bZaLJoT1pLPq1jvCCRWiP
dfuWw/YNi5DYAiRAZhZN94MvqGnVhX1jZLu5m8AcCtECtGDYLmaEAviQmX6EzJJz0MOOrKFHtG6X
l+PDIFMS0E1SC0Pm2iWcPuCZnFFneckWpvkshvOLhdxSKNRWfDxiWOo49pXOBg46sOP4h8oJKXUu
7MBfUb38wqY87HOeJLsRqGomyv8yt5CNQrkjTTUGWeCZWZV4g4AMEIb7lTPRBKIa7AVkBc4TAaCF
ZfBnBsm275DOdxPOM74kKvvNPey11UiXDmgznD4LWPjH8DCCMu5BONqhPuehH75Zfz/wK8PASpoM
jECvcYSc0+DvanyZIpvK6nRSm0QpQdg5/gweVUYef/9vmVgPz4w+Cfv8YvIaRYXrGdpJlbhDxHEO
uRYU21k9rq22nhULnp0PqzBgcTRpTrCAbkUnpvjWtAjTTwtPpePBcaz2SlysBci0B9RazKVhrAjQ
6UiaNGWEVhJdGQkIMYWLKdqC0UsWCMuc0MK+SOOnW+T9ef6sLFPnnDMNdRLexkPuGsVbHTygEtSK
+Jj904plW3lTUcabhmEXVjAoPKJe/Vy1CZ7s9q7HL0opAYRU06jdxuaf5PGsD4R1RcSJznxy4p0I
R8lwlpAICzuBJHH+9DTDbetEkR06EFYLHFKY9D3cRvukPiVwH2Rkw4aXAfKm28IrBtyAfgCO9HDh
8dIiyFLWF1qlGMQiQ5C3mKSLDjL70kqq3X61O4Flt3Hg7pVkDZiwmJohNvq9nfHY5gzWzWAqUqe7
LGZxX2R4fZrIU3VfxyAVYMFGHXKrzsdICxkFsYXWG+ViEMVodagmbws9efGkAX4AzmqnRSpcPDGF
CPCsGSyWCs2bAXLgwNCfsgXyrY6vVF3Oby1vH/3ve7qgHkZR+JLsTiHqvB8WKMUryt9xyn657Bil
p41amdKTuXeNZ3yuWTolSqpVGEvf+KtFACVeDCJpcQtbBIGdTxGLWIoqSXezEXKFS8h/bgSfkSdm
Mu4ONvEaOmFRfwojHnz21BRYxPhqALvH99nhs9OxKkvc59AYMRoma2nE/C1+eEPI9UH4kffou1Sp
OpWnBX5YBXRoim7PdYzpIKmnDzCfPlAwXW7VJdbXK3S83fmabEQkTg2I3OtOV/dfUWV943G+ApGr
FVWBseWet1CbhN7kDibG9HguHuyEByPMUQXtSL9OyIAVZoisBlG1GCvLyZ8Q0rXbVnS9Xp727MiA
muvOr+FznwZAf7NAg4t7DXYbhb3ByfBW8KPoIeZvUyP9G1jMGcElHYISb6a5zHv3MlYehMraSZX3
Nyok6vZMDBMT0TnRnDLB6KHRTvRNzz00gATIizjwCxsfjP7XSDdxWLN1VBk30ey4GpLydlnwsY8E
QMtoKujWqFIu3D08M/KEyCdKg4YWfOAlD5dC6cp20FzTBfLAJ5ajEruKnYUG7sFEjxEKjSCTsUr7
FkQsCkN/XPJNkekJEU6UcSXogluU7fiW+f44bfJ7JlIRJZJw7Af6oROOghXfHSBtg8WOqBMVgo3K
ltykBhmNVTTPyW2YEUSF3RhV9SEE8ybY0v9JKd0NKZKWduCiMQashkC9Cuj4UPGpDzm9i4cW/2vV
xjNhF7OlTQ9W5lp4V76t/qdiURYuLoAUZhEhrnxQj+QkXNCToybqLadRrSiVKyNeflAr8xyWBsef
/npZBElGTmmN9bJuR2vWMajFiwDYHy4/bdqvjSWyKvNJMmPO6pQaJo4tgXrORh7gxDc7uN757njQ
yxbMSmfnfT2avHYmYvJLuW6vIGSHUBQBiTqT9D8Edl6IK4Wj58NRJz62zEGHDHBVwcmflOrLmo4J
1TVP+JmCa3fLOBT1yk1h35PsBIiEK+lSGHl+OImYwQYk89llhw4E5HYwZKJhbqmh84KtpHQ0qY+K
cIwA6K9iSL7eALvQL98jd5ANuLHDSNV9hHjBnWfWfwOQozUmU5xLUnQbFK6g8bgHC1KPWbxXmbim
jCkhlubQPF14csjCvVqshEcAP5AYWJnLAHqoCwPJ11p3QfZAcsoWuD1QdN7ElWg5kmzFim2bkury
xZdgfWYF8PbURzn1/Vqck4HDmIKgJWP+rZNHckmaWlVwGoVaafhePVeG4AxNsI+VoP5ofGf50jqm
ynFHfXQzr5D5QvSaC3gq8tYcQ35O3huJW68Lh3LjR/RzoBWxO7dPXghctZvHXVP9t/ckxKqI7Hr0
NMCp7yCbRA6A14ZtMfPGKWsbn7XJQl/mfjl/TN/bHiBjYvaBsfI4DHkekiSIA7d0/Zzv1Yoxh0oh
24JPhG7IK5RKVWjw/WbPvPVnqbXIOoO4UD5twiMg6y5Js053NKQ7diNCjKvmAGRM0rc4p+xrX+Hl
isrSWVwUYLfaVQcj/pvzEaUy79xIp/aAij9LM900BFIonXiSvxLJtmprofMfoIqdAy7EkIlbiDnh
ofv52Dd3+qyC1Jfq7z1qnBWznhcmexKSbD0KF63YQPUErAfjR/dnasYWLiOEh2yZTu+nD2eIQ267
CqmZhVtitBlqXp5gC2JWm3zeaFgXvksL7vFnb6dCqamMeRSwt8Us9OjHItWhZKoJUkABYqWcgj57
zP8zOO6kRIqdqjocedmiBAm17+RZHLjZo8M6KSjGLHa587IcXbw62ZvRQ/Ftad7XrbjGhXvEMsUP
Wx6m9gaenpOD7USWkksufnOezFtad+ZnekF55GUtEDIqCC3CbYhnaynGJW7vvxU4gd3lmu+bFD4d
bViyHGIbMYD4QqijCmwlIiXJLA4xi6IYoGx411W7+XLJRGmBqNoQdOTzFtk5CU7a1BeBqjlZcqAp
2SQEJvAuuBWICQpu+9gQ93ErjVlpkkBpKiPcFuutWnCAx9GJjUEv+F8lWIamapmB9RrlKqJd0c1a
FryXRwohqijdM9yCPtusw3s2jPhUu84LeG7huKGdzWN6bZiJIC/W6KHHj3RtwrSbKih7Z29zmU/c
iigwoLzeIQwd9prCbTvgq0f46bbqKuG51eOBmLrs2dqZEAlaaV9hn3kz25Y8//xcymUC0Fr+l5xI
K2iDk4DKdhFmJNEuAimuiYu8ZhZuyUppNrpXcC7e7EbazLafvHUPEMvMU4LgKlB29aqPsMYPfpRN
yOyX9PAoW5nqAXhke4yhUogoXD3nekp8Qg84PCsKWiZNwFsBQvQ9HThHFrRdb+ZOqAGwO71k4++s
fSMk3+cy7WtW6wKS+3mRD2gSfK7gCkHzxDNHv+q0t0wGjHv53vtfmF1d9tG+Hgg7FD1ulD+3z4Sq
zAafjAwxyyBFhe4UShpiDo5ed9cibpzICsjx76Eb7TSX0m9TwlE43sVDjXV//0PQxI9/V7tPxrCj
mE7EHVrNSKZu0rFc0LbQwqcZCrwXxo/pPOl2BsxIu/1EqOyjq2HfjJFd5PsjMKWd2ig1bhx2NKKg
to2msKcgMZFgnittDBBb2gtwIMMdQHpPKISYug/LbnKoZfVqAi4fkuQ1mp4j8/Tjlgtq7g3Nkiy6
BD98r/LOeq0/3Tmx5HRsDq/9PzNFlb1BFLZ7gd1sF0oTH4FJNByhdGUUnPo1MOe5mR5LNsQiH44S
S+Te+i5TREfyFc+zTONnYRPYey9xqrvVkqwwZFLsGEqmRG0Yi/sMnCHP4U2LJzMLl6N0FUV5CjgM
9P5EYhjMoT256WlxeVqLOb4lKnSVfiEONY+n1aUhp7UZQ6wUU0JnLOnSSEWF86JAsUSXNpu1464i
r8JrsbIu7iZ7meypaDNiUPmKqcDzsuOoF1XZINCVJ73m/YMnq2LyYOEF9EjYUMPqX+Rja5RpS3Ph
qK7ljQpcnM2oU5Ie2/c57EGcvxbbBQ/3Zg1Xu2QHOssVquQ/FjvRQuj58Oo8ljcRGMpsc8r3Gl/C
fvgHC4R4/AKhpFbW4Ip3K/sXx7fk5mOu0NmNQNwoltkYeU84jt4V5VxXy8u5Zae8hgOvkfeOAGu1
2MlCoyvF2qZRujSTBVPP5YlVVmEatY2g4CnM+RtfbB4ofNCKyT4pUfkwmlpA9/p3VPrdVPGtMyOw
VSJ4XNJe3o4ryDHLV/+KKFOiY9vMTeo1EtWLgWDFs8sLd9M9w3KRig02Ml3HbYTCi+bmAVbKQPYo
Hkfim1tMG80R/fwF9ERQhsZEbuzwriPtV+pDPsyBtvscXjeREKDTJkaOS9k3F14EwPPhMcUZV+Hv
PuB58Wb15xDuKjsUTJDQFk/+LItmzx4KIoysAqTtArfXz2j14LZOkMO2EUK112kplBPFBa/WbfCj
A659PpOcEhs9tAXSSVXBDJWpUHVPHNJZ12cKohKtzK/MCYZig2TpGVUpQ8jnpfwLBh0aKQGDbAVu
r4MGwUE/ZQnfVxxE/gAzrQgEi3ATco2n0Kv8ZyxMvkfTYinsPDRZee0lI3Jah0unxOuajxjL+in9
sFR+ojKsWm/SFuJv8R5pWNUoC5PyPmhZ91fb2f1HdCgUIsbXUf1Tj2BrVVHXQcZGpKF8pRK4Y9wo
bFm0rvST/f1+92JqEMPyIM69d017BERTWBz6Wv2nOQXC7gpM4QS+8/2iHiaHEAuaFySqxxKxS5nY
CRroYIM6L8yBKQxpDIc9bO6wSva5B0OqBow35IngXjgK0ihMLh8yCMp9nxRhXApQXvB8IGXdQKuV
YgPMlTBhW3+EA9JsH82n4hkWPrHG0a5TYGCfPu5n0mypF0fvOc2iNbU21AN5FE/2tZuJS+0l54JY
ZNQEeTRYpjtHNeM5rDEf4veKrp8pn7GnxQKqH5L2QK5VJHmL5cIfsKkMPduW67dlid1jPvf2akld
aERVRJdJr4exgmYRFtRckx3Cr1YX5Btd71OACPL6WsWjjpP6TFPE3kLStKhJPaObOCsZpQFE1BrI
J0uxlesVbs8lNkmYOpLQxM2OevlHHRIiYrx/toqfKV2xxkXkdgq7JKgcd3LOiBZ/DKKRBQxdyKOd
vGNWu8fkxdnsu1MaT/mAp0kpDAGIrNx/dPLllolVF4qnGruSPIfHLA78sSwocxlis500EsYvmlh9
5iB3TxFfUPgiRwMpmhFXBPre0thEzHmf/fZQiQrADqtTZErwo8Jg1zfHoK03E8XdWtVLV64SKT1x
y4zIJsfSjaRAFRAblWbXsJgoDubOCndzqysY7VMpqlq+Hd0uByETYSUhTE+F2UW2JBHL/l83khT0
0Ry4kGVcT9YqIP6ou5YD2l5Dmxz/rR63Dqg/HLPS2j/k7rsUKTesMMivqfaZ6Bdu8Xt3KnD8Hsou
SrfyYSJqVDANCwZ1OlO7vErSrkg42PmFVb3wt00aeXeNASltY1JT2T5OEoXU6HpIXmIanKTpKjb7
8moRdOr0jEbTy8AbaC8xjHcRPNzOPNUQUuquaze6kHtHwQ50k2JsRaOXvwCZBpUWDuMGRzFGZ7Yc
MI5hrrdRz0im1q6b1JxnF2UJUuUIocHl9F6NZFUW6/ro4Ky4mbbANu+7oVK6tDkEFxYhAcijLG1c
VVJkvJKTUnqOOUbHA6N+yNgO3qOq8bG22guf+fsLXRmwNLC3zfT8alFNNdr2elJ+X5q0amhKEz0J
mCpgxoY3/3rJ5uT7al5v9UVlWdZ4aDK3Vz4z5TwCNSIVZMIjV9N7vg8DvRrXw+FV+Y5b8wfELmoJ
+vzBFkJFr4HWREOvnMkZTOUJBkq6YUteZNO6Br3mgHM0BtBQFkYK34PkmLDTUbH38Hz/27rP49X+
kzrvfCb9JvnsyhrehCATfiDNvPlJeS8Ymob9suP17DLMs5pgVod41NYrNY4GKbTXX3vQh/jhyTC3
TWk7VQww+rzUe8/T4nTDeBfEoIeLxwC6ochSKDJ078Ije0rCw6SW/eeh977qUOxqCw75xgCAzpVh
5dmGjXRSGgflQEal6+Zh4U5zUuASIRfRI0bbiDYCransOHH8tLuDKKgCgHrDZkzAtmgSPcCGeXvx
LR+X79Q4WmAlnMjoaSklUAYzK3EnuoFdCM2bOqYgiYD7qQpuTL3JFpZkfnXh/O6aoij3ursqKtlb
aEv2wn4noVGyWN6dqUHev/91zOY2iLTbWCxWSaYAvo7v2VdRMmvAIVjIn1Kg5lIAN70bz/nDDCAm
o1QGfGGPx6lMoFvQCJvePxkzSskCIQSXX3prRC92Fhkl91ZGJWYArYkCVHMR1nHYMFFN5yDzFYJj
JnQIv9eRYv6EmLK8HISlf6FSzfgoux8lrHGJH3IydZJk0zkUF2NrU86LVOgyDfpXFad00alj2MSe
aWWfJELYM7asLewiK0TSULkiXnQC3pZ0h494/+em0m5olcW/lzfzlyvLzXT7K7b9vc91yg8oYzhM
DZuvzGV4d0rzCsPJ3hfBmdDjr4cYMuLQXYXJ/n2EPTli199LvGSu/jhSxBOZ6VrrMlrgBbodUXWA
fE8eEK2EbBjpIMI01VXlQbxeNUuu08xjhyGmX4izvqLzCsexJsFh7Nq/QX7B14UwU8UrByQgHsg1
G0o/cLdksIK6lCuT9Eh8JjCzm1tGHqVpP7DtOHoZ/XkROAjFvV+1y0AvZ8JvEds7yyuRN+6ZLfzS
5WNfDarG4Y3Q5Wfk1ie+f3D7hHzkKToY8UtposT6dH3UEz127JjR3rc6yHBFqe9GGfy65IrLJoCF
xYpoZbR9MHCdWw5MWHWDc9lC7OAs2+7W8PzS0lFri1mxzzRBtfnUH4NmZSEvo18G+o5f97BgV5rh
klZ1a0SBGqAr25dRI3LZPL+V73JWAmSthiY67H00mQ6WLPKH9A3fOjEf5WCVFcTV93ifeIJz3pCE
Z+jKjMA74V7DYLU6l99/hnFoSt6br688t0qHXZVeIxuHICs3zeAuDT7q9aE8+z/CWMx0weeKrGmP
oNfUtDYNNaUpJjGgcgEeKMEUtP9S0TyJfOBHBmtzbenM5C+6pfAXWrDf45zarwGbn04QK3KDYqxU
S0UczyTMqsprob5C6LyGb+6tF/wYlweoqvAVMV78K/yGd/YCU6w9wZasQmH+pdWTol6bX8ZtmmBC
VAbVnnMhNFaO7CZ20xKfky2plaBYpspfYSN/Bl+GISoUPIA68srTqZIHWDqaAFCGtAo2HwSsFl1q
9lS8pB1pjN8M2YofYMoAK2kM8s6GIU/+520b+Fif4aQmHOvFrbdkF/fvGVLLwX/tsj9pQKd66iDa
2726NFD9ex/3832L4rG1+/nWhCKdnKSfIs9xfAbzcHMBFgrDaHcJAGJenXBGjlwe6oEl53lhvzRy
UtbEn1w/yPKQMNjV4YC35sGUSvUNbn8PUbT1o7AbHARRsgwj+366E4Op5WhqXU41vqUNOG8j4o9f
6c/IOfc6AFUjMcrE4MO9qqZnH/j8r0XcT05kK21AO7sPrO+DJAroOYGS9ZdDlSNkAgL97DMUveJl
hA6Q+Y5HOeX+YVGgmG/sUwqXuqXEjARmISjd7F1HD2qEdZSFE8OQnf2H5nmNtEaFVEE4ssMPpgeB
SAaNkwRFmJ8t2R5IGcF4nrjWuU9pkTFErRsSoBZTqqjso/WAvBbpuMUPfT1ZeyJoIi4xVkwF/LBN
P6GyPav9V6bxuv1scq1NrrCc9SeRNsciAWRQpDN9wWgt4D7CAKw1YQUtOhnuLL6uyXAgBMuFZG4Q
FkZVPXgmEldN0Lvm8nxGhYPkIZT9TzLPOM715KmazEyFdKloDOZNL2/wslqlIC+A66NMaFFmL/cq
XhtqcN/RApSM74RTZSubRwylAUiPcDJCSth7U9dncaMdct5ovJYPeOAVDgt55HWws2RA4E90Obia
TOJTTXb52ooGWw8b2i8UhVBaGDO3X05lCBh5wGlVbMcU3PTLxrEJuiFR89Fire94qLGUNH/XrX3p
qtF0EHG/a+lj3ykb2icRJ0neJbl+/SNRtLum1xvOPTudAxtE07xvLnF/qXmG+Ygi9nEgogg8DJD4
gU/5dz9QrHgTsQ2tlGStB3EDfrF9E9Fo3+tYNdNEuSYndZbEOUcAmfzQlB0cHWDtuCxc2NIbrW1D
+BdK+MtatcXPDL6DrQTsETwitdlRplxTVKvjs/2m9J/S6ssJ8nvpv+ykVP5ytl4ugzCfJFfs3HwC
74VTZgZYzqFtPw1/otlB55GOGAi4etw5ZJ4ezO/JpNWGUGGJ0BcTwYAEiLm67dL+iIWHWqr2rFYy
2n/ah6rYfTB/5qrKlQXEVqRDgtZa5mxbbCJSiIorwtEPrG+iM/OqogAK9pdPDf2Pw3Y2ggUt9Ty3
lQnvfWocreyj74uaVbwZfVLWiGfDCNvrDdEnD3l5yq04GzMlL8n8djve2ohT5SXxZxk57FaWshfQ
GEyWZtHnFnM+IcruFXS9a/v/C5Z6ZrJqC3WLJijyvth3Vd2G1W9qhfbkJpEB3AlSAJgVjG6fZwUN
uIY5NCsZxsWCaQI2+JNVfYfaWF9RCe5iF3NskIJ1Gvpypge2S2aGUmDBYZjuHZq6iZYsx/WDp+18
YPCHCgeAcK5HMA4EJgnn+FQmH70HRKJW2bxT6nlSsv0k8xxak1qB3FENFbO4q5VNI5ahlDCOKZsK
YFhqZFNcaIbtSti4zNscplKdIbi3s772zR4EiaFJ7bpqCoynLr2H0hvM2LrBQlp6QpkaQ1yo82qY
NFP0UObkm16HImtm+L8CUI9gmyWvgI7n9VsgKEi2bdTyTwcHu4mWMqmitWJ/zfQWrqUJL6+Gq7R9
h9QGwb/6nFLAXdhCMIf+L50JB88aBc3nG2RvrWNY285fNzywhvOMRqNIaozn65pfTh2w3Ws4E/pE
p2QlI1KA0owiM/mfBAu9wWetTIRu8oWxglyPJMZpiavZhOOTca4XaVqB87JOrWdRGA4c3Qm3J5Tt
PMeZltR6Kam7kyQNk9GBrCxDHwf8ISLXDHyucNNgARdYwGPM2XvQGxSIqGtpjhzBjTAkSQxS9jjG
/R3dk2f3IZLlHCBiysqQEEUvvQ0tSUIMfEsu29b0e8s4P4Apt3IUK8uWTtle13NWLJ1bKRPODVW1
t7d6c43JwPXjr9bEb5eqizd7NM2Lds8SArZYZ+ZWISiOEGYlQOvHJITaj8znknSe63VFV2piRbpv
jqO2nbQ0Fm2xMThuNq6wrgypwS0NiLMOKx2RpI5rhZvEmgkOMYzAERRBKSaPaWxEZD+Yq3WKB+zw
L4lk6aOmJJ6Wuq6YcfX2nS9elMO8u2VNJg9aeiwEbiuOM0+H7hpxsLePwqj0U2T6m4S/W7FAtuK1
VTlWJeU70l3q3TB41YfPn6gShqE/H8fo5jzmQLjpskfvGDhaEiSGn02cUQ+lIu0Z+sen66y9gtzN
xD5hTn+yEA3oNQaUiHmH4XZ4yZ9Mvuni0jWE+NANAdzgyRzjalmrz/IRB5/6BqHSdDALHBxVAmpc
YjMhNFD/8TXiXQOQuFhx27Fgz34xLhlAsS+jlNv9wx0+lS8js2xoASSMBfFxPirHfC31mrzrG8MF
DXp7gA+NCKkaF758jqsjTPwumO7sZ2Jhodj6G6Y2FM/RYaLoF6Gx9mWZd7RN6J7ZMGe4RSPm5cQk
zZUDjhE9wv5MXa6/3a/2OEjvNKsDrr1/Xam15CfkMDY3wReVrI8r+19zfNK1dcyv0kyYCNxlYJSe
kmsE6PoAt661LXUbF7gSdg2hnQET0yOIj9PmZTt8dW0AwPpxVhxzbTbZrbCM/xrV7Z6+eJvONNF3
SlccUDlZYcw3nOvxh+20J7pyw/CPM0MFpuVoWqff5WazJabtmDcfj+vVHtEyA5iA9+4tNdv+iYIt
dNPeSyLkX2VfFGHnGQy7CG+SycmJzo8CC9WJ1NMkMej6LtIfR3JMLyF4LXVKyPBa2h3Tl1RhX6ep
TRjSc8oK+NDS72Dp4tjupjyf8bMdGWJDWZmYHtdI1Pzu8TEi/9dl/4lcby8fjyQGmsFjYPXRf1a3
p2v41ryqLv1rxKbH66BlRFlhP3zhTVtadVLPb/Q5zZVtuDfTXA0Uld+FFmvNd9Y7i9R/NqpRAx1r
UUCwwTQndVstDR7FqEpePd8tp6RTJf1h+CRlg6sZE3KMjcK39ifJBjlWC/Gm5fN4qINse+UPSsbz
/mwTF2xQehs7MNt8J6vhdg4MGBULbWRr34kPOV5LwK+IuGH9TFAIvMopoNPjVv/z8/SXvTc9ep4Q
rLrWTzr5CWwJedmBLdMC7SYhw90fiWqRQlfO9fW5SmO6AreHwKeo+XOylSG7YvuqaQOTaqgz78Tk
9qzoiVY3C/oWjOWpdm9bq4qn412UlNRnRdiwE6EZRGOWCaNJcDGtacOHB4T5/4nbKxInZgailHQc
ScinpK6xvMZiVCMnoDohC/I20XFlAbh7giHtATa9uO2Jwa+MgqYMx4NjfhEGWMROkOD74MRYXa90
nYcECT85KL/sDDubXMPx0tsICCIu5ZePyHvUjdixJtMX3ENqLXUxrVNxcdjgjDYJlOpNTZGtpBah
P3qhHSTGsIpFvBEARrqsHAM4khLW2LBGXr3O2JneYeGh2EYz8j+nHlyokOdp4wJHAOcP1QbI5Z/2
pdyl0HDNJQqboj8snXs7xON+cj5jrw+053QOZmPQV3OD7WPpKyTXpZ/d98BxJeC15I68lVregL3y
s94oaStf1Eji5FP21039QmzW7ve+C1bpJUu1ujBMYR/go+J4nk01kE6gSN0UUtnRQ99ffCxiShJY
PaCiPNiI5fOy3dkDI43a7wmsDzqLIXq/Mv4U2HHdBvELRwFf6IPBoQTzviQv2gyKHH+F2d+LlOgb
+e3ncW2SbAHB3+JR+PkvkbOF0XZAir6W71XcYHs7sR7NDW86K6NZSMPg0/PbxJnASCSb5Fomlw1G
/TvesFkG1z4XHrDK+TDV98W2VYXokYYTZmXRoogNpWAYP4nsmd1Tj8w03uruumIHUbk32nNtxNvp
lngpGzPCAOpYPp6gGNxxGe0TYvhQ/Ip8mN9AG76pW96YzAuRNR5o09WznfzUyw4aBSPaul5FZbHv
rl2wqII2yVoSAy0PxmxDHusyty04miHakmv9lxRc4kH/YuCgpIIRl/oXUl5ib2CPTuebhecELXpA
oLSNwa7QwbuPCaP96ZqAEVtj7/X53d1r53K3c6nsnDP1qvqLE0VbZxzGNg2KVdMkeEmlaN9m2V3+
JCVRnj2opmESh0RXwEkxmWoYiocSdNA9cQhEF5mybUVID4salY+8MYSUc8Z3/CuO+OsTbKu6AwFl
I/C2wQIszBEbcqS4FPjLAqNPZD4QKTG/MpuYINZfI3HRufBBdrjQngxzrdk6NkUKCC8PdJucaquE
45RZcikjAoR+Bsjf3fZcx2Nc2oY2KAcOODh1JMkgxd2D0fIQd3WPl0DGJlLnq82ep13ZZM51aFMg
7yMOsHK+Bh8fI92fstVcvOEcnS1PcFXbIhpL7qXNtJ7Pty7uU9kQz3GYx33Oa+GZ8MvOQkpvp6UH
JjRDtgGFRyjpYKABE2DKBZRzGJuUgBTOP3X+obSe/iCFs6fCBEeHDs84Lme1BPI1R7JWIT72ITWc
HosPFDi/S6aIwvWuTaFVyjSaP9yx3Pxh+ckGl0/a4CnwVHIG2xY1/LvRRwwDgXpZmB+CV4e2FBGN
ixzd+kO4LhB+ZW+/boE9J7S94cbMLhCFp5pyJWys32y7MwcRWxW//5aP4JuynS/rQd8HjRItJHKX
6tdq91T9i8uVAYGMQliBU9/W4Qk6nLRJEBxaaP8phBFZK2mxVFUHCUpvGJ4vgl+puZ1eoQgpwC7w
H8mofb6Cw9t8Zl4aVKKwmMFR17ZjoiePnh9R9vtB09RQGbuQZXoA4AiGUAsWDMdxHV8O49UksvUF
MN7sdgjcecY2LOTfJ/Br/BwSHtA07PE1lehLQCMRnTt2+JDcLXyg8fxcwmE+AdfbFUkCDvu+L4uV
C+2uqZSrGKGQcW7fqRJWRXmR8sHw4zpRQ8oFklUrTR2CmvtkDEUDTTdB/gBC0RLDozkpKhN9P7Mq
BGejZP3rRetTsq8S5IQ2Pd13PwwiqgEWfK37+b0A3H5OmYvbyT1H4zPLki0xC0UF15Fd2B5J/qUM
ihLRSNNWsLvsqtTkynu8+LdHdwDDZcqJ2+KhonJAQoDEqVETeUbRiuy37QkLWJWfsqNO0ob1NtAV
phqMOSc9CLQBZ1N2W9ANE4sNDbMiuWjp1Zoe1zjaCHfkpsYHKeSC5Sj4OFYtbvbX9e9D/gH/iXm7
mPMOjhX+Rcx9IxcgMX6gazK/Tdlx629bTqLuW+Dms+hG0JHnZ2eaSf5D7GKpqzDf/Qwq2/DK8Cy7
uEzFYVeiCT3b1v8ZZAvhJsAP+jom6DECjheixzoQMvD7JYkMCHiROfoFBSvVWaPMZ9NHHCJmccch
EutoQ+GWnniNIQj7z/REFqf5CABCO3ly+31e7XVEZpesBL8bJxZXA8FGuHFA82/C7h5s2kc5OZ0s
ZvLDFFCQlrIbqb/eCtkJ4psmgh/ZMB9NXs9taWYiCuxlm9yJGs2RqKEOyfXGYryRbzSNVlqnijIu
UK40FSJeLnakFCKIMr20Y1k1UfkJd+KVEEtjDbtuI6UgzMCe4pD56/ALBjcz7XqFJHys6BXU2cMy
D796+UAZ28yWzWLAAy7ZD+5LkSpz5MWIQHqpXPT38ImGwFr9ojUdYS4eXE++AuTT3R0sC+ym7cfm
7CrhYJ0HXfP32quRmKUM0QYiEpYbEowzhcUcRjOPO+bPEBT/ravBDnoVW0tAgPMq6wVu6sAAEWj+
qJHr/G5VWe1wS/TrglkiEdUhePld3QYSD+EGX7bjS0Szu1a/c0Jpc1V36pVnXAuveNNchvdGNWeZ
xSp312zigBUoHURQm1I9VEWPty3mhlN+MgLNlD1eMqUv47Cdn6QcWiki4oO+0/FN+4rGFKo6YOr/
hEBrezx1xv97rcp07xnkwfLLMYj1tIFNo9ULDnE+dBeqfVnlHvguoBO+Dwu/eFcY5ck4ZQn5pANw
SB6pUjGz3SBLNF1CEHUPV4UtvlynyZ/g1J1Yj28FjLqAJbFYaadqLjXoBxRHSmIXKP0Zh6fJYs3C
akxGC7GH2lrom2CrmDOU/dIpxrLPlfUvHMUZNptye2lxoBkFu4kAGpcxgctBiaX5e885WYKU4odU
HLNwTru5XPCSZqhsQmxk9xTLDDuk0fBBXAPk5K5cT5gWSIh2v6Isqmx7UkMm3Jy7uKNR7Cn2iiG5
Rn+5t7+n6IXQ+VVaYraLIWhIpzwTieVsZ8c/YiRY/XyIvHn6XYuUhGbnjeSYmGTXkRwjeZSzXVLH
Cad8jdJVJz+yQrqNdLk9HHmvm7k75LnQEsmgmCcybsgVbTRkB1ukYAm3xisPISyikFJVOH50aSEv
hPEJIsR+wvGPKV9wn2HVjSoojTzecEflKTsrc8L9wqVJnzqv73TKB9PuhI+FFoRqhUIe9GfOKg/6
5UuxbC9rOgQA/rwQkn+cumcklO0j6ZuDKmxQ4duZh/DFsqXKN+RcmW3hzWFYzxaw8Fe92Fl0S7qa
1SAjOKD5xabgZD3mHOUhIrqn4iAST/YeutUmv1+N+ZjQmfD88Bi40evtJQeuRSh4HHvZSgHQDKOo
+Oz1uao5/uwPPA0dHekO8QAVm6jBZA0vsn3difwSrjZqZldZlGI/z58svhgQoTnN7zPmjXwCAhxl
pocCqZccl90FpArkzn1i8igDpmQK+pWSLrb3v73GZADLFHB4xCjAPdMxp8N5wNsF+7HEmHEaVexw
N+LV/hHD/DpL9dKRXESxAUY04py9YPrUKvpVNXxMnfjUTg1gmjHyzGDACPA0V5NKMtkrLKUtJYvj
asrLkvBuR7oVFAjM2QgRp+1ByjUY7AOlCG7zcXJaxXn02BnU1BdXpf6wb1WCi0lj/NyBhqsHgG4H
zc9XJaHN+BXC+1B9ZSW79f+fCAp8AYUz+Zhxh9pbg6S5GdxAeOHwn+WMx/+vbrlxtsb+MgIuS0Ht
pZjS6o7mZJoIWj5bZsPF2PMd7kkpTQlu54G9UeWvZs4wFCDmwk1wpVF3DKpJGB7oT0bBoE4F//nu
YFre6Tt9gHlWylLH8wolAmE6gVd66/GNqqvMdC/MlVPKM2qJGBmeegnvqvo5glcFIcEZesHTNfFC
pIAp3JIL7c2FNAriKd4vJ6TUB2nsUKLUXn0LfwLvLob9wFBfsHGsSV6ZooDfKibFT8tSOG3bWubu
hBzEeXotT75bI4X+z0lQcW8ISYQ95qxk5oqBsDXwLvAnK+U6FmMIZQ+CjetgFSEeaaeY906TXoUN
le34Jpz5nxHlOy477fDTFdv44X7TMOIF1PyL0cYaABK1MGbj7ETaXn8QSyi6uG8uCKjGgO59ibfa
n9BY3Q9l6onAHUGe98mThHk/wMM62Br748ICRoJyOa+NlgDM7sGdgg1+Acv22s07DGjn4xsQx/bx
5k799Az9h4bTE697tVDavWVp2YttwmeTMfKRyGRO0vw9bGkicZkxYtnu3O7hYkVHSr9VNS6TItfa
FpnOGb88I6BggVdI0/wDHP1hsh/Am1RBpptpPmtSF+QTtjA4fJteeqF00HqDV50ub7zN1GFBGiIT
XXLG24U2lu7SD7fnoMw1Aefv6bqn4PE+6mFZ+WqhPQn8N13oZlmrLaH4vCQ3WUiqOUjxLVlyewYG
M9eaEk6Fts0A3DXOxzqGUbxmoqJAOvOj5e5BKid8ztPg4ypZvRevdfrJWUOkmIYx8e/oO7zXQHBl
2IEEk8eLXcBoZRrhpIe6A2R8yGN1WRjbi6sQwLZI1Bme52eT2TaURMp85THBwQB1Iz111/14Soha
ITZq+S9iE5INGRBT1bOY9/W7AsZ+QW4yXgPDQCEexDOuNV9gGbjJu41ezmREGLilXZ8pTCqivYBx
hI7KLyIIicJr/JlkqSPYPWpfBe6GnHmz6kWD5ng1ILj9j8cWNxp5HnP4APGW1E0emn+GdrmIuqdc
8NS0Kl+ln26Cl4OGRC1BKZHRqZ3YqmDv/ZsdDMbw30N7pIoBOilcRY2llyMSFVvcW0Z/3XNpXY/G
0l9skgNW50h7QQy8dOBOJ15c6P2Q5X5tR1DO9CWGjSmBV3xuMLuhNfDGBS0M0Z3IrU92Ov9jeQfr
nZnb7/PEwD79vAwPhO/fBdjUmdDaZBZUO1qf8hPg2wxfDFJ7w4y9cJqzpxcxHaQCq98FqYqAC2Ui
qHKpKIBDRhnJeGTsyYgTUcwdK3eO8RGqzczsOMs7E9sP6AGytO0w4YBLoiQPtI5Z4LsN+7srIelv
2yFXmvpYacUJ5I4IVA+Tv5hcSQxGc1mmeNgq+azWeEwVUvJHG1hc7a/Y3Wchf6sj1fpCy4Fj2NRF
yHP0Q+9m4g7bCirK26HXgrTatstVAChXyZJS6Mp0iHG8d/xqfeN1vfK9zbVy7bXwhGtDbAY+t27d
01OarhZohr/U7ZXs1k4o8DLzEWMAhSG4hJBwQz9eyR0kyFxWV2PBDNUjgIV2a9gltu048qNkPLu/
1n8boL4Sf8Zb1HhOj9X3/aHZ+NiVkyY+LV52CAVSQsrAIgQS6ajOgusTInvjYMARaVmoCVqvpa4p
y2CytK8TZWMivyzhqSpEEI+WU8N/mYi/SQDuUcD478hOQqsw3P4Vp3lEoMgJlevaOyJZiA2toNqN
1AYgHQ4zBfVe1qJdX+7eUStJdxepsctD75h4Kf+U1z/I6mD6kH1BbEwJ+vTZEOHs5D2PUdNgs5Zf
yqLNLN6tk62uo+tfJ+KJG+ieT+R+YD2Zr7MmbDBdbMZF989Sd2eqT0DE91DF/3/jYtWAfk93mLq+
vs1XBv3IQ5hnDl54Zl5TtmzoF8Gxm0hviw8Ktwvr9xVWpl3LA4NWiHo436wQXghT9m02BJe6C/Uc
vfbNr/SgtSdfdLQKJ27Dqfi9yEDkXfr2dYN2hez5XHzsWHxpbtHMCvhxPMu0y80UFWxncdV9GyMg
hqpFUC7AlbakWEx7zdlk9EGsn5Eps92Di0KEMPBvnZdAvgrnAFffBesu30/oZev8jSXr7HEWJjoV
O90m7WWVCd+zpNAfTfDZ68Kh+fkcTXwzwsKbg/PZoqS1NvZhHXE7iz3NbUVcXgXAkAnT0LYN2u8L
bajlo0NJ/j6NzQfT02pqtj1/pAgD7kedmSjWSvAbAqlglmkj2ZwcZYWJKqTAc7oCh9Fj/DshVbQc
V3cZ7C+psrsUEmBHIDgLNB+0basq5us5rjpYNJYifkS5svNo2/Y2WAD3IPVRMVOrtn1m0pAfRd4A
QcGJ4Uqgg+qD7MfVnhksqatRPpVw2v/F9l1OCDqSr2KgFePclLG4AUaUY7HezJPi/mhb6Zzfuz6X
2WXFhiQINYFBwGVjadiIE8X293wIzshZluAPg9JtODq3m/XusrF1JcGvLmtpt2BeSPHazjkzNLFA
fx6VIKhFwH54mxzlKd9TTV/J5A71qMEXWyustVPQwVcxPKGIYEVCSCwqCcoi3WjYkD1+3vKn2NUM
cAoPjhtlQ9WyhjfURV1vWk6cVvG+322ysnk3/Wfq3ZLGqghPpXeHMYp4GzFWPyaqa0AmP3PmCkbh
UJrMuptBP3ZTuGzdfppCoZGXoPy6veKMIbU4B6ftnvc4jwbAn85wPc0p1miltJNtzrS5kjJTHU2v
KEsabbobl5PrBYUaD77XmaKyXdttwO1f+wgSZ+ylPqGPEWCqoEFcSJ6jtr0hz7RYtTDvn46UZjGf
PnltnYlM8XF2RrMR7MXZDbI2hWJLR/b66/hLbp2TgnCjyU4MbqCbmSaosBe0T5AAAPGXdYW+j8Xi
RRdRej+k47B3Cg4wKuhFsPfbphwEWy7wITImRJ+UkkkvIco4lQhd5mijIyZZNL9r5SrGV0uEhhOl
Bv26dsBFB9UdBIR1CfnuRy42OEiloWHthLm09fsYp1ZivyeNqsj+D0K+o/ZD9O7upMhJq6BNQ/Yd
uKn4oC2yVB1gOiUNdNAkOLJzOzvPROb+aGGBQiYbiXrqggzW0KRjBlBBOimdShfjkIE+SUuc7oZD
SleLl206mSUp880uYLYpfTpht19Tv0eYRswyxKhDTGtL+WTOJwqQrwJzPr+DKEvmfwvJK6R37vrC
85dkHUfyydtwBZWR3QIJspMVeUZ8P2LZXGiXGNY4eN8nympZltcH2HvBussHgbJFodUBhYye5dtA
B2v4rACT+28jszaL7SKyJPD5M1/LyvoZQ2lf9RI1Q0wMoQquQliO2TGmeBPAIdubf452hqO99rjr
/b2c/UCxGpbtmZRwcCOOKjQRL/Ca3gNKQXJq4GdeoCp+0bGlSCHGv1wJri+DozHpoTYAUbOStja6
ZekfqaloO85xb1VdxAWAjXTCeZkV/OYdznrr6i+7VXooaJkTHTkJYL61mp9oMx26hC/dLHxNrlRp
tMFLvJs/pxI2HK02/qflCb+2shcnUVg6QCmhA/QZ+Tki/5dTDXj23lTDkS+nkiZLkNFFDQR3PQSH
FkvkW7ynreNzbDp4D7hIvetOamj3Mu8FkE3R6E8bAaLq7rqJzJqX3crpN32FWiOlWlI10fwkK0PG
I5YhhfAxUC3320Wu7BfN5GDVsVKWqxmnPzg/s9SFdRw8A0iP4ZJ+lcfO4yD7a8WSZ3bnG6spYXnW
RkHVbinJd8qA0ymZuwmDT0oanH7eiuE92DZSIbIu4RAOcLlu0yp+UQrRUz7LPztjpmXN/6kSM5Q5
MsoxOWXw9lmvUVZGcLNynXGcHyiNVLbFEo8daVSrxO9oEGTiMl+mIgrBTaStnq1WH1VcoVlmrT7f
5rXW3QVu6SWZsIP4cPyJIeuxjF9TSh8jleyRMOdItRvewNHPjSgX518yGb7X4T3AF3n0aPcZwJyH
soJkGGYVQwPuivWplZvLxir+ZV9Jb+VsYsfVXIUT8RXguCAyf6kOhmp0ZyYwwN/wUS2h8mv3abwC
yCpEsnBE2GuIY1jZW9BnJJItTGGKcUPIxm8hy8MDJym+yiOoM23YAC4EsHA+8k9GCUVe6uSzcf94
zvuiO4OeJLJvvSbYfmCuOvY961ro1oi5ZlD3kejf4eG3LAHIjJC9tjv//W06Q+1e23EIEbZKbWe3
5SkLPbYJDjYS2NKzu22Sb/nKzC7m3OWhUYaB//u2IF/euWldp0i8uN36/Rx1T2nrh/v5+ZI3qW6I
vas6EcxDnl15QNWE2bxOyDFDiA2waumlBSMc0tIwxvKsNnHvgyACQAdcTa/k0HE4+YZYpCAtQaYq
EaIbk0XLoMNw+z+xBMH1wsXsOgajeGf1ofRxsce7bHaw3h9ia+a8YntrvQ3tWG8x9xhJIz/VzJWf
7+RqP3iqIkmlUDhyXisteQrskf58QluQuuHyI0uNm/4b7JrB7qG9imb44bIyTdRolYexgNvuvYiM
X8Hr04OXckAsNQu4tW6Li1e1CCP4ctf238msX3xf77fPs1LyBet9S+Z8a+5Hku34vatdK6THW/vm
FvZpXmMZ25F9znzvyUb+7co1CyaSyZtoEFsZMb8/8oEm7Ydr1u+82+USImwIjieqZ1nnr75Kctww
D+dtreDbLpKATP5glnlPzOnGetf9NBHanR1Ysyp4X4ixOqU/QXV4iMXmmvbpudyfaOwoVmapl4Hn
3rckIQq4K4y/9w+wV+Jxlqk0qBh2UKBTtkP+aUSa/XsXXAKKPQz4BYr4f55Iu6pvgDYwIZ/8C8mz
5Lw9JHnHZAWpZ8jtGLTWuv3gysiqjAeMJJWqKcOOmJwU8hM3l7NWkcqzdikWC7tEZfvRpopRDpFL
NRTkKJwIjOhnL0VKH/fC8m08yo0wXPyiPpoGMQPwTVJtBT+rtEwfA3N9b7bql2ucp2riehKwRSK9
DUUOmq4vjA3g9ZGPWzmDiPbr674Sq8qk4UQwIrIL8d6SULW12w8v1xw4dch1z64q5Y29zs74nABB
3KQgfotA932mcj7MLShz0XJ4OcKNd5yZXYVhKZIrijyMaqJw+w63sUT2TLsS17noxOzV/ZarIiia
s1YkTsewSsdHd5EPIPrpSBgs8DN2FEyPE4csVTv+zyRYgdIuQUbgdpfQDFqiu+UM3yQ6H4ioLpnI
n8ogvWTYuLXHCOyJ6uvxlB8u2OfJ1YlRq6Bm22sOiYtR4NAskcfSY4X8pbolWhaLgyBPtt3ajri1
IcvJy2s3IrG9i7mkWLJ3s4NkMX1roHkvokTDLkGI2rODah/tUjtsuw1PMT7fJ8+AueCwfRn4p7qC
BsTi9Pns2gl28zF/bqhnjftYt2eG7nq9llNUU746KDzOxx53FfJr2rIX3yHxvsY0lqlai5BDpjYv
TOPNPzjzaFFJ9EOZ2gKyMs4WdgA8o6Bz76S+kh+qZ9+rMA6wicl1SDD9LmtZqdBirLX+KG8l/R/o
EhcuRioiXLct9KSAHHBT3oR0m+CdnZapN9SPZxSMCcnT0CS3gE2pz7TS5utKYxWjUBbj0aQIsXd0
axdC0BoNbZJM/bkY4ak3X8ApbAwBxFouSR+OEM9fr+VVirTDxc1EJkR9AgCFvxFe9WV/oB0FLUtU
31BFmrzet931YGUWxO51NeRO2LCEvsoYUYNy8U3i4FyZkEm4RnYw/Xi3t4ZkWP/K2teZ+mpy/qng
fEvY1Fxrp8Aq8SoLwaVk/HCnOsSWeBy/i3UP/6n+9gJuk+UWAhRtZdFv4aalusOsxz5ant+Dmhc6
7MnaWyIkm6B/45nph1emGuaVz/AnXbo/7pk+EEjKVsT8oTycfR8b5fESfWwoS0MW/EQy5lP/72yz
9BRP2+84LOfhfHCbe6NCxO43mtGunEdAeGSf39GgSf9jChJWYqUTXBrmkPX1ypBIMhX09PeaPHer
apRJhPW16/AGu27ZBnFMyHv4+S//EbRVjmz8/4QNpjO4+BeWzPrbM2XNizV7mRLnj+/7K/xg1eqn
q3VR1YF0o6D7c8rfJELleLn+RkNEbFu20LYj4X092KNmX9fkUO29SLXJlZThi8297J0E00FULPHK
T6c4flPEjpDa4SWSib7FrIrM95/jFE/CCaaO3XXPysKHN18U2JVx22DqH5tLs5PKJr1Hqf0G+pmA
6CBlNrv8/cjXbKg7k0fYBmCey1+zBHKC92bsRlxwUpVMVRBAkp0zAZYv3GJpTR+ZD4Cr8u4KPJR0
rBZDnfwcwc39SP47ZQb9VYlbSaF0aV2eJvVzUhW7m9S8r9khEXbmtERliz+PrgQGD7JoRjDgoCl8
c1HMdRjtMOgzBMa1gaSF5dPOCwuZpE4K7l5weJ2MuxzEOOweJllTMOaYf4hx4/VlpjuFXr1clC0K
cEHglbV6g8DmIx3fgbwmNMFHCPczWnuz5i7otNcurzG9mSBTA2z2gw7cwd9Paw2QSNzwv2uM16Jy
NAgTdvO/kBHywePdcDllI6pFTHWk6P3tZ4fHPWAjTy9LbY6zgKtUR/YtsXOavcXgjjcySiNKkjXH
8Dird79cxZM4zTKiVLbkmDPjz6ZjScBeASGAxQmjhEefbvtR1igTqo+JEMDLCXh2p/qqVgy/YPkR
T8HC98q8Ic99/iRcOpxARGMSGhTAfxbLYX4Fj/5N0hCfzBs1EMqpQre7X+hboOnM7Z6rNajs7Ebc
biUabx7DCLMWrgIRT4K2KTsyLAs7l9+OVUkmZfHjaJrIteFgXtQ+dmKG5D4ks8/JADp1FoNHfBSU
wXx2L/MZxOamVKxNZwbCcFF+/sS8ijKjnNNnv7ByAOeyxfPuHM/wKx64Ahuy5l7QDJDhYChhnSbd
Dzu083CFWqKm1Kx+Ymo+8Lf9Oy75YtrtEGkcNQorP6NHdPLrJoV/y2Uv7aXtkvO0iLWq6dUMA9dz
/jI6U/2LXRhpL08x2qPlWBWOqHietzh6IoTFUTo5kAJUuLMRAdoud5KkbHEkEbYqvUBeOWoAe/LG
VH72liye09j2G+eCZsuVwP30f0Rx5tVp1rdCYBSS58HGtzi5fXudtKQlaeS2pl9HcOXub/SDPjVl
IzZEbQybm0fbvblLIdUn8CPt6v8wG5YgGRzCzbvVxgkuGDY1aHy3WBmsWjWjRW/GEVKmc8eSi8jD
+E3zV2MN/+i0JXY/RXIuUVIAKYdKKvjxjX+tW62ojx+bNL/VSpfLq2IFDzZpcWrTp9KXQyFRxDms
iRyR9FxyvxkiKd45xvkbiL6Ja/Unq5/tAizh0Vcdn/81AanbxNi0czhgkFKfyy0iK4pVtaLS7NUY
vDnVg+hGFXuMdE6y0zwWE9T2n1pMeO3sjn2OBq3nVuMC30MaH2+SDbA4KfxeHUOUXACzciZ9zP1v
5v7xM8IXIguZkF7fcmqYVHUvphX6ZeW6pZYz719v9e0B510aiR1yR2XBKGj/5Atvv9fdtTWiCPxo
43/YgMdEF9Z31Nl11puuEvhQBwyYcTgV5jO0/qR91DJiStZoaIbX0Bv9gwKdwFsTcye8fJlm1ewH
w5lu62aaBs/t+NWUmNKJuBjm87TXX4npnE8Bgs5FPv7bOdhc/iS7I2LSucR7i7Oph3q5WBQeYvy/
KO5YURs2hQE1h2+peYzo4Ji2sTai1JbRYKfxywLbxS4Zsx1XG8ckob9kMorWLyP7unV/j/jAwWem
cgfHD0UHEIsLR/62100EjXwGutm4x29484yYLKx5eDhh2wHIAT0jzIBapSlUqqy+nPbAA97m8BRn
/YDNA9RYMqKrn6bknh+KVS/jNDGWfAKA5ZIgaZlYYtAyt+6/iiKGsmdLKCrxBpZ75/LAhFT/25+X
NFgCrmY8V1/Fon9eRaTyOMzV4gJ4czPQeLawyrKJDhkDidwyvrqyCoVgVo+c6qpIzDUpp8r1w6k+
saxzyRHF1bz9llkzQR/wffrnixeSHtNdEZ+H0duakVLT3I77nSTNROgobnMp77nRtwJ+h60eV6Ry
0A8rW+kMnTTJvTypgKj8vv/4/o8OluXBtBbBO9SUEnt5YR3oJRUkxqiOnkuToJPHIAOb0Gcz1H6a
xKwmb4+aMGzu3WQ+lmKCOhSa2T8yf6h6dhRTNBXIezuhAygkVY2UJWzga9e34/85BI9KZ9ZcqRg5
coWzJP7ld9glSeyotFUobnrILvfSkouErzAklA6NHKVYWrsnDW9peurBQSg+toInfuK9WIH506z4
5t7/YmxTHHG+tjGscLGeZ1i/9QKlgEJLJs8yf+P40uf4z8BY5ESKQjq3ir+VaC12mhnng5ceRkHY
r0hZ47Neco6vF5Sw3ZZ371/dTq3Ax4uU4MSQj7NUUg5B1px5VLzN6Gl++mYW8YTIia7xneJZ0X5t
UtFHPvVp1p+mO1AHZkvrMkArHDs0DDJXBfAW9cOuy5wZNfua2arkZEXT0Xr+sZ9BxisTC7hxDyGx
Nk8S+2kQR9XYUr1W+qc7dJLAME5XuJll/OiX0OrBRyXsErCN1KoormEjauj17syvSkNz+5WS2zc1
gWtgDMjkDAbWz7tzXQRRG90DoBPm7iV1UtlhaX35V5s+glgUIUFOZ+14ZAfeRTIFYwX6AVRjXeCB
zfIRuQLLNfaI0XLyfmh/EPLsuPuuUHVgF9SxXMP4ZONG2T51l5AVT7Z3sVXg2BBkWWfrqocBnc1K
R8a6G2KLAEsEzkjX5KZ7u8Jahv5qgy+F9FeK/IYD73tgK3nTAR9pIxhT2LQNN2XvIboWDx2OohNl
/sYYzSeipdfZl64o8Y3jhu9zc61HLaMJSNIWKsvM0z4mPV8+h5vqe9w3fQgWM9FA7MTPlJSE8869
ttNaheRXWG2j0GcpOdy2SnL0Gg/oX9Q25XeI8NIDrLI7K6+DvkRZTsnK2BJYllJNVuGHjaDrRM78
fr/+YZxVcT/Ix5rWdwpAxxxWxkv05loWCEAZDIrZJafkIGOHiYAnCcBYhOnQT5PHEu/Mc28cJ6Gm
pT02uVrp/OHxQlfGrxP4avldl5tRyuEdTAI4710/N/dd0zSNXVh+CLRYuUoOELl6But7a9V41dCK
+ESzwlt3d4R+M1GdtO8F9moZjjJqq8BWPP/GROnRPynAfaJ+cE6ggUMdX6x1ZAki3nOO/PYqhbif
mU++q86+4qY0Cf5xV2Fmye5BGd4+WqKlEI6Ow93rtgFGkyTeaY/myx/mHl9YY1Dt9DOoeanNShjV
vmDZ5U4+s43UVa7teUH7fvuCmJlCn85hGt+8akR8HKacCrQKM5o45dFNPbL0EcOqj8AUfYrpA2jt
wQ1kbC1buj4CnDEseb1FAic4imYNl7pTIykYbUi1rsA4HEPEzFrFjt73gGmW4/DFLT2LwvOtYVPB
Z8tJQkoEcf7h5f9BjBiG6R/0B6djBOJvIpks7a26VfRLnvUuPMcuY9ayuPOL+PPS/Hf6RByZKRFc
GVbpzmAj/3Q9YTSjeVwgRuYQ65/PpYQcAsDBwUTCcrpKSLVJAaNfYyqVmb2WrR/6uNGUJQLIAT/d
qrGkPjNqE8Z515HGmVqhP4df/6ubtVSE6tq6ILc2QOy4ci/NXbT+j/K33wPNx3lk1sEJvKIemx/z
dn8+dK3jCzJmnwoxum2aqxhiom8d66ftoOMpnOqyMquOT93ydPnFnSxcx6lFYqdDDc4JlJLr25fX
EZjHjQXCRPdvEMkAsBv3gJ7k3oM/CuPRX+sirM8cuX+k9ey6oE8KPWUF70U1fIzAfGrXkQN18wIX
r/mIetc/3NgdPeNKB9lZosizAhIuTM+RWLOi+7xGi1jhN1YRbkEr7MkWWWndivvJf+FVjR/nv2KC
5mpbJ7p7H7oeVH/WN3wItTFW8iR5HoIRvBrua17FpM/Rt6MtSsjXq3WaCbPtxLxwVZJn/o61tGku
pqPEvufyCHIvV9bAa3em3Mj4K03Uv95Q9DqRvdXoM6MVbI250YiVd2VlUobr5ANr9BbBOnPXmP5Z
suATvj70qKS2vRt3jlF7MDxfcY/IGVBZpeAvzJ9TFIZR6TYkhlXuKvSy2VNjupEQDtz65cXS5B0c
V3UywVeafGGMdiPv39Hmy5VOD3mHVlBdd0lkLueuYjtnwVyEh9eBCuAyi4Pr+BLBaIvfPD2tyMYm
Crqruzvl33EcNKjzCGlgE1uHiYlPDZu2o1SIa78kBqW+nnVKFnjTjw5LZojt07igMNF8VnfPwtFv
zNTb+Ee7BmaAT4xpgiQdEMH0y4mfjAsQ/OfIVCG0P76dt4ROwazidNC0aSvtgXcM/kIZwkVmDMoG
eKHe9duBblHaCAcBsQDsL1RqWusRZxCnrI4SatfmLD8pDqZCRyPNbz6/dG+q6uF5Hoav/jJeC/no
a+r0K4BVykuZ+HjQDyqdqn9NV0j7/oRg3NGE4+beK3NmXXYJdwtsc9zCHEmLtL42szKY9C5w0aGV
pYwLMOP2Yk1GBcimUczx/kGTj/qq1tq7o3cyS7PBGttGgldVzBI4IIv+92I5nBuavtFljsEsbVMO
m87i8aPWVMYjGQ/Z0TalnAZapRM2t6U7b2GbSQ6ssXxn7Es+OMTXT8UUbf9cqo9ctGpT5OTXQ3Sj
+kLugC9JjgOO66KodWUqkYzbYuVoWV3uuQgF6bA8+/DkiNICwOx39fjcuy5xrbbZMhK71Stk3Hjy
QvLXvqo3HvsUqynb8MbweS+biWPGMiqnb/gZhfu8dN9pX0mmSJ3aiwGzEvnLYBzCep8v/fWUY5Yf
Sy9zNvuW+ZJiHvTbAd+wyQFQF5b1KkKi1JH+lgmEQcWxqbj6MT5vsT5UsZz9kbMFCpp2KB1IA8Sc
rm+VoNF6AxC5VKNsT3gp/lmzoZggdAdHr3sPrVsgjcJcm9Y5bRtHDi5z24Eh5a0R7qKy36fD6uCF
cPWHO1sIqVL0tCrTv/krkGdQ9XolAp4at3ayHK5yf5Momqms/anfoN5WGmq4t5WcHkPVZal+PJv3
i2VlJBxCgrXXBSoP0OPpRwLkrz0nvkzdnN5Rf5iJ52Mm82o23xw08RSDRFKbXZl2NjZ8Dmjo8f1d
Es24BPgkzEu8cXiemtMmRH+hVBZx4UXj6eIEWZkeaMA29SZV/qBo1O/8v4+lyRgqRboGiZVLnEF7
uLsbZGuC/FxO3UUXgvBkZZnrT9migPBd0AIAf2He7MmIvfIG1aL/D/EoIOCJU1uclypgn5j+Zep2
CsVkkquRg4C8CBaqvY2pu7Sy/SIG0a4PP2iVLRSH+Aa2hu/D5D7fsvc4bnZHmYrN3Lw3QNNV0oID
6cggN9QQtzaqz/FEVklnGz27NAhjjYsuWuUp2twVZsqTmnln/O70M8sky7dl4jSDZLdFMPGnlFMq
JDVFixCz9C63bGrdZc0t2EbFgbRE2++fSlLYIzMBTrYy1NonyhS26598oMHYgDVljnBOxlfWazFb
K1mpCSmKz518GEDZyCup9VTXy9cC+CqY6eQwO/R2zEy0Bg9LnFeLauj4aGbNiSM/ZaBmehqPFkSX
ZSukdr9f1rrm/wpQFzLrms2649PUAuzIAhxOp71YpEpF45lo4JT7QBwVqRCk2z+C8Nwd+zEC3nxx
RC5jJtaxV6MS472nlHFJFNp+qhPkWXcwUIL3rpxG/JOP935qBE8Ple9agZbOjV5QZJ/8mrgeMgbz
6EbDXMbs2B9ld1vtUwDhPvSTCYRyQz7xwbuKbc3QaKe0b9GE0opp8xXA3QzZQyH2WV3FfyoR0T4W
oThEiVDw+4+U4OZyPHwUzFWPUuJGVdWXQU6Qse0G47rlGuH91QgXvqFhstt4UBxbCrCWcMczkVQm
+q1stKhoLH0fQX2ooNKjX+FGP4jvF8xHHO5fbaxTkiH02vGFqnnTaVttWXd/NRMij0qH+w9qsg04
GlebJdG0iDM6FIiGDwpx6jnv1jdjdzXSBypO7lEzKxFfWvZcSUzELUB+V9ukSCP/2NIxrvZkcGDA
hkKY7IHp3E25n6OMiMrhYZl34iMWYl7etMRj0HSIWcPH9zv6uj7alUXGxDjFssNBiHySBwR/sus+
Z5wLWmQT1NVrroHVAvRA+BLlDzQ4cQo6vWH34WGCgO0wTE/71RuIWVdpTnzUMDb76xoOui/zyUL5
PohTuEodzKN5LQOSm4zD1vSzMoxD1IJ+r1x38fvsjvNxfm5pTrL5apW11d2IEL3YOWVqT3zlRLSf
3W81e7qrXyQVkpIF/Us4yvrOOSWESdY59OYZtpLjauR//UwPUv7KtRZ0HycJ8hJoLLEOgE+IuBEi
PQ1k1YgQCgYz0wf2EWJeSVuPN2yVm6dzABUR76Bkln7sixs75LfN6FXNnCvprx4Ik5Z4ZsrVFZgD
aqyzfJPezkmMRLuwJhHtk54OK199RwSTKIjjSp2E44lktunJdsBtN4p7WrSKc8rljAZgPMaOKvRX
DMVsrE3+dGYkLBGTzUDao/tKWCH8LG/c6VUh451X5BEIqgXLAgdab0dUT141YN8Gl2bVOUryX7QV
ofTENS/9DJfgLx4qHqAfAzlmAkIPiWkLhUbMHv9XY0CvB9ot9ol3fnz/NU4wtO57c5j1dEoILC3C
cUFTuZpHAFzlgWauPNe5nUdRwxkl6FPzLvt1UIkArfyCE1zClLgetH6eW4vLg2vCmrh+3pPlyMkt
svq970dNeu57LjPFc7m1U4/I5Y1ITm9ssqN6wY5nXfZhZ2eE2A/KU05rWhmA+9eAYQDrPuDp3OV2
QY1ETuLSAHit0h+XCge3PMH8iORsIf90+UQixRGohmeUrmPsaSB006GQnHSQM8CmI+ajQt88XaB2
xlF2nN5a6A4ULlWigwEKfHAanNUq7JA41iDRGR0e6XPViAi8gmChnYS9TUO+dPW7gh6A9iSXI8gj
9AhU/nvTxghcJq4N+dDQMYx+6s9FEw4UsdfcpBg0E2tj5Kudd6rI+HkFbxHPko2qmNx/HqqodDrH
ZJUc0WXo1pbWhD29tholNe6o4hiZFuTLRoD9YLtsp4jAG+QSY4n5V+AVVh2RI/9Uev5V+jZ/j5Vo
rUZpH9bzMbQ+7h2DXyWhmu3HMRgsGh8EVLDJH4lMUIjTs+5ucnNyum+AviNic8VKLDpnHxnXIMMD
89Rbl+cGFz3GZXDQwppH+tp+UgFD644/O8ZqFogUleBAdJbS3SRBDnhV/2sIzYi6Ds8kqCVc0jka
RWj2eRe5GJFJMrLL6kMfIEIhy9ebOvhZG7ysDLAfJPJrGvUaamW98L8sjJDvLxZdD17N0VVbxbWn
1/P/vM8wKOYzXmAf1mq+XwI0nXJ4H9mbtBnJmjrDd9Ae6RkKlR8hLOBE+HJwxGTqvLrt9XSUug99
MqFw0CJ/aeaqwprN/400Yt3JJEvkkC7+ZUtYJhREUtLC/E8XWPKQA5XJZJxBPkZYQNX24W4UIbSd
grbzjdGsDvpT5IQDBxmPM2Y6368+LFarMmLtJsqszKR8BuEY3ar+7k5QIsDa8FaeaeZjjrZSlHgj
KwLxnvEadULOHjOGGvb303cDFJv5PSndU35u4Lhb52tOUeVxEOfAfGfY/DfJosXluyua+xIY32t8
dbVKxdtzkZvVhEQJRODZOFvNaiT2gZO4eCivb3FKnJpf16WS+k4YrCG3J1zWNW/TIiv4OHQuN7ej
rLy9zcH5Z1fhc6pVMkFDpZx+hD4BxxGcLcDjGS3fQJP3M+XALDo+gVXOfWLC8P8tk65d8z7Vl8eb
cTTaqLMFoQCaEtKXB1pgLdTWohsPlsmJmWIxAcrAb5diWnx3L2ipx7MN2vMWJ0cfMoRd+2zcrqZS
mqw7bPRJQ4D0AfgrMfxuBOt/NyJKc5Rqmx2eCLbqd1JaL5pXLgNaC2hyySzzgbWy8U9j89NLTzpo
rnvoPmR2q3deN2fXFMTpEay0Txpi0mafAApBd+nO/h4eOx+k1534M1i1JAt68KJwy8EbQz+XdVnG
Le8L1kAbMLPGrztKlbCddGjruk9QzyGusbYNE/kW//+AFnksa4spCipR4GiazHcqzJ+tg800reAz
6S8zDZ1/EADa/2w7ciJRBgxfiYz9xwEEn3e6Ut/3qOBB2ObBVQaLYTXOSqMhYeudl1LecoHeCNx4
FQfdTBKOlBG1HRidsnxP04nI/sxLBRTsjhYzBw2FnKRJsocB+jpBgIW0fozdhhwsC1+id3KHAInl
mTQmStfFeRMgpKORdotmfSJLGvQNlYHk1UC9uTJ+ry5JZg5MwQIMbqSofY9/YXioKi+SmWX+gLqJ
f6S97MbyV6aAvkseaXBON6BlNj8pw0kzyM8y3cgA8rFMn3fE25aV9LKQOggCoroph634jxizTF8h
cIk55TapEFlNy8cVMuGw3X3camKJKQAfWPpzQsjwpubacfsNsOSpyDS5nrTdhaE/MlLZrMfmqIw3
8454BZTov0WInmqDDTZikLRPcdb5hM74FJ2O9zAY164Cd99KoDI6Rf5Wj4ZZflfJZD0xxbq3Sgp2
y/bQjmwaZUBxYepMadUhbqHCsltG0eobWi82XZzVyP4d9nEX/BJH0s0ka5DriXto9qR1Ue+yeVdE
o+HIjaG+pVLZ/uS6ynoPLaA1TqbOd+YwF3lXp7MY6XyISAQADNLCkeNk0/0WeLlGHQ6g9kedgiCU
Qgel2Mt1f+A/OHqos6SAyNJw5Dbz6cG1/Sj8M/HECc8zO5Dqzg0OS/8wR3rZTyG8clfvylyUF/PW
sdImsIToBy9M2Mdd9GPqnIfWX0hrhWKAqQksMBWwWNGdiCvYNZyLCf1uDefLG7cWWg5GwI8uaawZ
LSftDhvsTjvnb+c26HyB4qbCldRkSrh2H0M/MihYybQkGLmjciRHtYrDl4p8rQO/S59NPMW25I6G
2dOGuEP7ile8tdFQKmWTmvg1k0D0bhczEJQ8djZEMdHkKE8MN5dKyMipfoFU0w0t6y0Ndm+0XCnW
8TIIiZ5o2G3Xm7CCxjNOJZLU2na3sAnmuu6btYLBWL55qDUYPPRlyqxl9+9NH/z+6BpJcfraZZVJ
WjxcOz2v+ei/9tArweoz6b7e/8vJnIvCaNmKq2dHxW/zG2kPXvGgEHPMtgQo7A9f5jPtIG03hpAX
gjc3fitkOfOi6OK1Lp3En3V7wXoQjPvKhXKOaiJmdfY5uG/hBehaf2zYtCpoFinV570nAXOCHUHx
hNto6D8p9illEW/G1kD3A9WDQo07I2ZOma5fvWnllf924PyIbcqXxFcY4GFyrclI0uH18OvZvtmN
7grN/mq69+3rXnjC+UtkF/vNN5MKtbNIjumihDvPwoGGF6mLyDG1CyVnqfxD2XHQgBmpRxK194yD
RejGbL9PtjOHDcFtj0J4NmELt0CCtNtGiIlSflYd0YVBMJdmYn6Rr26sZ4um8gQrYb4BrGSe9McI
8ZgbiiCcrel//MOhi/ZNxxLXIXItJSD87N2coC8khKKSncmDW7QNT2/btsxw8CmIgqEpwmkNrA9Y
GpIigmrjlTpWiOYYtHyxj/NnnVes4AxEv30I9h22g4QdKfa7+gEHx8t3I8Mh6ibvAyCMsVIZgHBs
kle6qf+gcfYOO4SegP5arAx8nL5xo0cNbKLyI4w7UA+kVqE3EczEu+EXef8XSNA+Tya+CIWak2Gz
M++XUZaWKnBhcituqFQjMXMVwgjzd60pTd+Mf860H22lan7zsWtV0rqWG+kpEDnGlUp7fmbbT/BQ
3XfMNS66W9YJO4GX9E7NThDiGSCjK1ZGfzeZlMmloDB8aEr3dmPX1Pk2DAFMo0Rs1MLEcNiKmrUt
hFZMDsZkDvE1CuwTVsbjzDcCAPse0iUjUHDJvI82KvKYTmogi55dRjLw5DUKeC1uEhze12Urul90
CnVHnc2C5hR7j+vmA50hOLVJt22YQTtB+48Cz6XoaEufmWIYtwXa+p5gAg7ddzBD1itw6HLz5/af
zK9Pu2vzAcXVRXCR9Mh9SQUFKVL5KcLAnnuG9v/sm2xPTfC6PQQwV55uilqBlT7rAEhW2YkMkYMF
LA61yO1MeUln0it61nJ4LADVFt9NmjvDARKg7jt3BYyKlW0E9aQUdH5t5QVgFra1RCWLyy5uvoDL
LZ7tBIwyuSt44RWRdd4e06lDDO7BrOUM8JoUviduU7PuZx0BI1919jCBPfeB7EYfdG7g4ldbxRfl
pd02iaLDNW7+h2UWVmYu5vUPVBmDlFTnQnc9s35rKHrbgfbZa0SYgc3q1j0Unhn5GfVmBLJoGtsk
dTdJz8wNz8NEhUwtnOPczaw9uFI1WO48OUR2goYJh3LXr9KMh+0QUpplS7UAEKUZ6DQyQF6YNC6m
1ymkOqePNIllFGoYqRDuj8F5q9UJuXmTqy+eIEjkz1PD3YhhG+zHRuDyiJLhaqbyjh18kCEjJj5K
fj9LrmBMLyWvZeLS1aYt1AcOynOZ3LJk1A8zFIcDA8zprP+y9g1GObk1TK+3SUTs0lnk6+LhoKMn
QD86rxZYoPENeYMJ9lMI3WyG3RXfaXMsWgxmVWHhiEE/LvYK2pNlEnZEyAqtb0HQHXJqkYFcWu7A
RYp7gRZNxuQ8x/EqmMj2uU1J+U4wQnxSUc7BJE2Ge8LyCUt7AlRqBDUftKJ3M215Xz/ltVDpyKMd
wiJHBderLXz7PM8bJaE7s7pu2r3F38voQMKFUzRGIJyGqMLaPPga/t1yIlBc7YiBric0xQnSXhCt
yEMYZnGD+CMOpEEM6wDTtql1QeywN8IV2Cm5+iAt7EJlUhqaQWv8ePXgl7FNlL13x3cPEhY7B632
Xnq8SIed5in8UWd7eyIcOMvXWwdZGLbe+hixorEBvXxDFEO8WDOnwMZFbvFrVWn7JaolDlmiTeOV
SvydD63lwOWErsN5Q9vZMRE/0bLWKmK+vPN8cVYrXq2Ad/JgfUvdtkHwpVwKaQ7jC+qV0IqqI0MT
zGHfLkkrAWu4GVGnoFf5x8mnbUEE8BHQ7FOgzBJUMQ2TKrs0XkJaetxEwJxXE51XiuboPlMsgZWN
cnDuzwvjKKONvVJlDiTB4L8UQvoa2i6a4NAwPy+KQeB+Qp5OjTf8faD4b97cRWEmo6AS5DbEkFXj
NLb22fqB1frFBIpggCbBJX10iV9JBzot32Q3EPs9hZh5jibUigqfHUNGnuaTA4+pR8BaSoPSx0at
4HA8V1kQH9W+67EWh2IJVdpwv8gw5UmX4IFaovoKzH4DBB+S92EKkkylWtKtzGWmgY5OA0KcTo8i
7ATKEzTDzCMdVi9hBNplG0CD2BXDBV3ru7KDLlryLRE7SZCE1TlAzs0Zp0ToDw6x7JfiHAypew/1
UltG4/GJUyOMc9ZAqirFUKBGOVpkQ8HZrFqR0JqhTWl7jy6J0xEqBlUZ+jYHoA515M2jQhgSttNe
WqHttjvWYFM8TqkJQLY+6hv0ousXAXlGs2/3bVpiqL55eDGf0d6WGfa3gA5S8EvM07kym65hQXCd
kH6B+kwRfaDHq2TNV95ZdtrkJ9f2vyLFRbUsaUu9gvCibucPn1P9scXCNlI4p9bRU65XZe4ByYZZ
r5odR+xCCZQ7hanlv0unlPz8Q8p0Z5ZCqBkX9g5M21z61y79g/j16SXiZ5t9lg/1AF+WX3eZD3D7
kE9Vw9goKOK/YQryeUwIm7QdtwK25UOU0pKgyvvdIBlbs6CVbIWU3becVpj8jXAyq9L5J+Yj0zSA
NPSuSY41BapA1OMir3uCMFnZVxp45aRj7JcybJT0VeUfrfXreJQsd8BRn8SMi7aa9FTg8guetBG0
Efw+Ufe8nGksH03vJlC4VWHU4ERs/gpHQXBPzltlcdMbWU1yVbfAEFophiFu3XB9UPNU16KdRkoC
BvEQrn7ZgS0aVNzFvJJsldQXih+xqTWoU3yQyDmEUHBZfyLUVuTLVQ0Z2HRqwcnhSMF3457elWYV
dL5Dz+RNiMcyEi2nnLtaOTYWRFPed8XAOUo8RnNplhmE8R4kMVCLc2zM9JkrKyOLnQ1Ox5ZrayCz
xs30T+/3h1R7wyPjAiRDcMSVizFNo4o1IAbXotgztQFvG1m7TrKyE/LvtXriZHeMYlWGq7tR9eUl
OkDfi5DJVPxTaizFELldEvhemn/5sREInZcLRMcti3P8912zBuzlbjBk/Xd/DKCGkxEzBy0vJHUG
CQ2rASfh0J100bmf96PHpIHDC9y035dmLawOMXfcO9xPUxsqmMvkPo2fsG9WY6Jo1OosJvR8dY+2
ZmdbzVPTSbQdKuE35JlokskqUANnf8GWygExRYk3ckyH3LtoS5x34IKv9tGVzsmKflcKbyJ7tIJl
BoZ28pPRLHH23g0tr1u8ugP4Dm0co+wM3etoxCpfyWlnKTUainCZQZe95yE6DUZCst0TzwjZFapo
X09SwwGV80ChWRqHN65hZV8q8NOG6go9et7U1hyf19woQVX7mX+4UGyourMKS3YHgBKDL8rLYAqk
H53ftEq1DL4FO/ho4pBkVS5tIvDc8ncufqJgzV4NZFOsNtTa5TdNog/lLF8/94Jb3lbGbW2I7M1T
csgy6rTvzANrGUL5iPB/L5HBiR5AIlM5rKg0k4bfnXV0Opa2peVh4i0TMPZHycURvFkSzIWyL/7d
6enAzLa6inzJktIs6ACHmoid50r4XWQOEf+I4ntHKEYfAQI47C5A+9N9PanMEIpSbwL8Do9rarW7
4eaN+b0lC48cgMxq/zZHr0gEw2JMnJK5vbxVBj2ezNAhqi3vsVB2KeU8md27DKdCuQoQ8nI6FwJi
pEVVdRqzHgI3rffrpO1xzrtvyRL58tEPsrlN9evYagxLdf1yqtIyX9pKhbj2EKZ5+7nm+6jEuhhO
7Srz23l7ZeXIA/66HwWjU3FAtcPqaCo49zrWO292UQmPMB0T6F2TSXbFVWa1qBTTETCEFAzojV49
/wiaM2T4IItijVzn+GVNWodER5BrayqFP9NwIScMD7jvrMgjvi1djavuzsoyuFQjkHec2+Kj9wut
jf3QCaZy5DSiM6Vfmb9xWc/TOp8dTQT6zU42JOXxJj/PIfqDBZ46gl9m+KDMlzVd72UL7uk+fr9L
l9tRqhawI6n8g+d8xhHJ3CkGUaaAtxivc5qekrv+bWRRQEqQcQ7vEhqM9Y+hZwSRs1K8AX4/0njD
2ggAWAEXLe2N3EzKGa70XbS8b91lSFVhcvYwy7cW2t2HPNZZrUVlti/uhvGuNnx+XLRf6gzYLkcG
eXXqrxKmkmsUWlXMP+S8snKrCvp8W+ygDV7KzGe1myC+j/9j2JaAlynAhSJ1TrxiQQRdujTK6asJ
+3qZLZgXXCS7UVcUSMwt9NpWHlJaR3Yd6pLwrvRi/nOKMyqcYZPbg1USO7azVHHzZYBAR1lVN/v2
W+V8wxeDUB5ntHzr8KKDIullr6OLTsepwW4tHGjkolrnR4QysIFjucEv8+Q/tKjaoBgY7luHpSpz
BaqokKGUaELKFxnldR5j0xXs4wzO06a33arkOSyr80Z8Cz3StI0BRxmPXMSc0VmWcCyjNSQ0Fklf
e5nkR1lz0O+89UY92LI3oPFyFcQPYAdrkInnao0UhfmtJ+8C7gzy8IGiOh8sUjDSyye2DjH1zGsp
XWHlDaF2lhqnLp3u25Dd12truOcne1A4N/OCEz+47Iefu0JqsGeySwDbJ7uueAzfW1Ma2yv+rezS
3dUV665ofulsjG8HUw5yLRm5N5ZP3clJsLeEJ4pINPYfUEuHxFCLN06YExQwjdTfstuaxD2EoOuW
LaigfAOt4YzrCMDls4T95wxrJQlmV7rGsRfpSatY+yImcCft1dXIv34gvOJZcS2rVndgVlTHdA9d
1HHfwTkmZ7IWnTz867O+gtY82k+iQRvP8uND1QLT6hDt0+qBGijw1RFhzs4DSXvhiZ0k3jIv+Kt9
IgX6MOMR11+Ao6brTb3yEsMEc0QlX3pGvRR4b/JAHos/0FCjwhe9AYP4OcBrmyMt3Gwww69cnGo3
MXCFV01zjPTbSoJHfd4OzJzqJDrHxMGop8YnspsWazM3iYI8mqQZ/WfR+T6AniHu0Sc2WTdVabER
0pYPQwEICXoc2tTg4TEghcNY/CQQRDo/ZeJWqxGhkiAuiiCz7NqizfXlK5YU260vyeGv2kW0HSVY
Oz0fu3VHj6LdqXm1s7DpQBoo1Q2zZdibOkTs8Y3HbYvquoJJaG+qHaMZNFE0vPa8I/x7vWxvY71R
T5s33EmGP5ImhV1JGErgDE8DHN5BMRPijcLqqvnAuRp5A0yprqr8/MtoQYbxjPjOM57rBx5NXTA+
OoJqmhJmaxzXJu0s/QFRWlNZoDbO9bXkz5trfrd6X2yC14ppACOte9BAtHbWrwmUqKkQpimc/We7
e3WI+0+R9cb++CcD4/IU9MXYQnbWUQC3VJqob/TMaXv0B8sHtz90SRHDxtKCAzCnQUm5+7RZe9R5
Qs/tCIsAap5ugU7imqYb3DbpjztDsuXwRoxvEwSYHqREVLifl5ewKBnVsRZl3J0kqkVy6EiTtqfN
HuHBYKLh3VSkg8g7sieWRkYyn9U6GdeDDMpZhRLFGWOkJ1Rt6cVRs5TM+5buKgj1vWJUoW/9Wbc0
hYx2XwE7RFn6g+gcDgRRC9SCNKyvAEx290Iz0og9X4wDqW7s+TvBHBP9So0Gm+nqSglwesnSj+Nw
XlViTEZB2EEs5M9l9bNFGgs87RtofNOylpBZ8HieBL+Nd/0MysqqoZSDyXIUIxKKQzlPLTKcCzem
GdUM3yWF906AzM0848VhiwSWZMCv3Lux1Au0fhjlAc8XoA44HlhVLHtHohiMRyZe/Lzm+JtbabFs
r/qrDDJFaAvMuKbcPZbcr/lcDWgNzPcEZlZuKOM5SkujEKbJ19WRENxdnkXsMJ/ZjUU3V9a/6MaZ
ihMJmPOJ1o0TQwuuQ6DzEEurnyRetBUbIgXeF3tDk6CAlpGpWAmJ7LE/E4eqrot7zJVtyB/Y27Qe
+vm5hMyPjubRvbPRD0C9SAQKj9Cplul9aCbjNrlYY2+nXC/jJ78qLgMTnTXpe2zTisp0Yq8nCVF8
4lypxlCv0JuPRPL/USzMzyWu83ZI67uuO23kItWe+JZptq//+ih7ORaDWG+TEP5MuuvNFS/VUvRh
5DeGBMcceFDwFLQdYfZljjnk/ccQWgFXimAsMvCCBFfsCl52tBDFqQcj2Z/Fmcx647Zmkro6iX0A
PmK6NI1jdK9yVsfCteSvI7+RxVxt3FrN7+WcF26PZrCBjrR+BxFL0ojyyxjko7S3a8qjjTAfsQBT
lLNSFXsNH8q2gnTAl7uh+qRkuFU2Vl2cGY4cLf5MAwDbEfI8DkNQI/zkUzyHEC6USip69VdgRspT
RVEnkVFSp6ZtyyDQPoqfoZCy82rWM50MFLQvU+V0U59sRx5RDf/WqDHMgDDpH5c9kHRUUy1LpTXf
EfDSJyU96Ro0+Q45duhGaTS68I7aeozpqCs+c3RcuOyHWZuyh0BT4DBBHlROhDXY2ttVA/HbgCuB
AsXJrA1wIW7ARePPNGHbt+fMr8VL7bmF5cScOjfObyAKIuFcmA9KrrSLYdtYrRLQNnPtUlg7ChDA
ubDOHoyGwmaf2Xn4b2PNCGyst7/Qt+9EAnmpgD/qOW7t4PG4JQCR6gna5ZD1shBbhPTkEfbHKAN2
6m0b2IgydIlk7axRaK7YvOoH9hgw7tf6mz+BttZfCMKDvK2HaF/tSGMfYbVVUa2bDfy+xsCKRG3A
uHI7psXVxHQLRGUS6sRnwt9xa0eiy0gCJJyM7YuEmVZF7h0Te3zGyxZ7J1b6cl6oiDPQeUmf86dE
gmvw7wXb2JVxbWl5RoEU2IaKbpBIX24B+wKk2LFDnx8UWzpq+usP5dE8UeGKpLocmEErwJ1AAFic
0fmK0wj2Li/TBdacpwtG0RCFbvG2Mbczsbgy6k+0+q0TWdTtNLZprcEFrcbcVLfyxjYZ2g0oQl4y
py2mCbOknMdRVGzlRoDJ1zWKNO+65HWsaQWRgUnsdnS9DjTMhsrNq+I8bftQ48/EioNLsJpKTuX1
OjDghxnR4uiBF2S6Ga0Qg2MYkqhE1aiQMand6WPb01GvD4graallcvn8kQBXoD3tc38B85nj7Kc6
T7X0nsninBT1JiNX77wEf1vZysQGr7X6zO5C7UsSlqIw5svwVMPew3rI72pKuxmiOgiyft48iPja
SZLUTwyqxCReWdSH7RUrl9K0ipQx63ZJAjIcmW9Epkn/sBdVul/fNJjSIjYy6Tmysih4aOiRlQpL
ZgXOjo6qfGjzS3LIoZ/1fLqlDVcqWEIF4VQGhHv6URGeCHoUCrg9BTw1E6dVEhnz0B2MHGDLRTEL
6ecnXOTtzTZMSmPp1p6zqvkRlnbHb8dpSjFvPs6cX2sZe/2904oa3nPRGJ5kbKeXBu84OjlwGPg6
+fhHy47SrBujueFWRtG+MPhHUZtcYFYK4uM/BvSS36dO8YGECBuYjz6sT0pjVFmGVBelV7bYCu7/
uf4KFTOZT/e5P2+fGjAelMSecbRsIWULXGi/TD8gpMZ4dGeb94LcxlTJX7cTjQW2RpKK0/A26M0l
PrbaPANaEg5HlM1MzEsBnPmLklroC+7I7W+IqXZxHafXbzOL+9nBBxAlvUIaZZ1EMQD/Mgt3p4qB
mCRck/MfFwBW/b+RY6ahQgc/8ZIk33WwgcT3MRPLOcKvlvN05BYPujCCVIoySKQV+YNmoSAI90Bv
K78GCcYnzDIucZvQYCAu4ZVOqFsTdvb+6FqlWM0bSs8iIM5eUdT+6CE+u3f73e2sVA7Z7m0xMrdl
KBQoiUMKC3qWXaO9tQJwjeqAq3FD5KkogzU3sFZAhY2lqu27Vu9FIZ0ft/jEloAxHy1adDtfbgEY
GDldQ0vlJRQtHfWIo+KEn661xUwtU3mzauMMuO6jGSBZQJe3hw/FvSe7+s7a6EjRdgPAimcVOhek
a8gr4sQax66rfQVZtiO0fbxVk8Rw4PvIpyMUuN7xsbzov+9iT3mX2C7XvTBjf2aVmSBYpwGpmIuB
67Plk/FQ5uHW0HsYH+8Ghyh03lE5jFI1WYi03+x3/8/AlvS1UhrxJI7O4qrbuG3zzNq2J/ZWjT53
qTmrdg2i1PLCj1SVK/pG/mLlLa4iqxIMGseLxvXWaVYz7wXbvOtTQFPgDN47vvkl4HiO8wPcSAPC
1NrZjx5zc6IWCZuYofUEth6zcpmJA4Ao0GWtFv8F3HYpzXiGgtjKpx/zi+wcXWWthTSlwRX788yv
/yS/QKmOftNMRXsaXpqexXNHRIeLh7CxwHQFLeON9jJkPqK70K57n2s6bC8Oc7Ae9KnAeSjyy8sB
Da/XnC97WVEfK3qx0kiLz9rw0ThULmn+GPuNuR4EPv2gi7disSp50VKAaf3mKSUUNwx7n0hIoJta
XQrmdM/8lf4hevkSPD6vHXZPTLtindBDM8K67n8YirqQAg7HAtDKHNL8rxo6S0JH86vcJYGQnIm7
dLJGocEKzYkpK16G6jA5Dmflvyw/DrWiF5Gfz3EpQMI+hDFC1v0kcrVfszng0Vg+Lprt1XnQQczS
XR56OJGCj50wrdEmiEgk0s2hBxuYijuu6aYpsyjbskxUGXOetb+6iRW4VCMVfm424525K/2kpDrV
TTajyPyhtnQLLDtaaTH5kQ2ULC9gGGr0oQs9+PllJueFSuuAuQU0+2iWFsIJXsgN/hd18wseXS2V
WRMBMiAwfLUYpXGRFLUEkG0Q0KBnyXV8sGshS7Iv27NbXN8fNoPQJYMty7t/TdIncH1giGSqZ3Jl
ZCyx+4PI6QbhdlA/a6D+7k6T5OCAqG2Zd5hL86Xz9tl8TVeuZrh54Iuy4bO1XZM6rj9Xiz4hEJC/
U1V4AhIAvEOhlhbsWgORprCPxVT1ZRqmtIvzhQl2iW/vkBRJIEuzJIfVm4vmTli7zBm747TOJ+L+
KKp8Pzyb0zSSMKb+jJLbERW8lb0n9+5Y0ozN6x/de2R5giujC3QejO2MQhdXfPC3+A1/rc7UXBrV
T8i6kFZoU+7A7Ql6ivwGfj4SfIRauw9OoSbZuSv6YUIpSNcEUlNUlL4Z35FTm2oeFfG9DfwrXrY1
ZANTk8c68umz2kQYm2HeiCfU9wFkcLxLNTwbWuqywQFwf/Iil8KF8PpGzS7OcejFh7A9OwYWWEwf
2sexoRc7RMTthPQLXnHjYfTadSkGnScJvjqERmOk0ej9a6hlPasya2LYXfvUIlf6CI22tqLh+hK0
JUIQke10fiXbJLgbPdTOw7RUZVmhbGmTLUgpMQc1cc+sSVk0iOQpv78YXwwvAJHXA0p1Exmi1M58
/6YQDbiaPB06qSp4wEg2ZWOl3FXijeLfT0G+p82cpaZVMB5JJYQrQzuCUR8Jx/diRk8cNaYN5s8N
Hqm3YNleWgr+p7dge7pIWKOJfhhPqp5IpuHGwerFqYf6ZF9ilctgAP6H1b1Zn0p0rKlTUN1bKW6b
YmuPfvs=
`protect end_protected
