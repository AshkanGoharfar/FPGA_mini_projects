`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
ZBBntvzBw91yFP/qsR39VxnuPuLucGFMl3/rW9o/Y406GP0GW0tCDmSKDo6N9wgd2bpu0lKGMhsy
j/vmKPisXQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
cxTph+85xE8haGkAAbuDkRChhZlwB+F8NeLenEtrDqas83FAij/meDKy86L2nYa7NjC0ANSLLLHc
HGpR15xnDVXQZIKxwG0SPtseq5L2jKOmqKtQ6e6NBhip9Yy+ZIv6VM/AiFNrMSHz7g0KRquL9YRp
eDxmtp6JJtg0D3bWl+E=

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
MLqqfGT7x7b4jKea0bW+SUI9aIyjz1K60o8IMnDLnldzr6DVulYxf6Wb/8a4Xnk0ej1ufRVx8+6u
ZUaRwftSv0Fbsppua8pf4LNsIGA4mayKOyXyuPV2JuFKGjUL38iMtZZCzTNeD4LejDoLj1BI0dmg
FhHJwhDV7xA02q7zHjM=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pLxdlMySVG8N0wmXk1ZM8Ely5tMuuQ8upxYCL8i9Yc7hYGpi2MsZ+a2Vikcpr6UneNIX+pcOCB4E
PJfJZVDdFbLhldW1SIuWRoaU79CllgyGsb0TMpxZmNJvd6yXgs9Z7+IJVuwLgvEukR36gTzIAUWR
yqzJVbK8xvCukiLOtZ7SwxjWbp+IGwmT9O9v0pg2jMZF8I/zfZHrnxweNvDk11H+Xfe8BRtuJhL+
DBdy2SCbdHMv9CbzUSx/Rt+1T0bi4D0YerdK7iE3Radnecevs4fjs1OJaEIKT7gqkU5eA98jeNEk
NDYpMfKZjyUV82Mp3v+OjY1xj2L1+2GW1ORRjQ==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
bsTximibIhmxUy03Gl6ANqJzXjyik+dvNaMC2SSO8kFuAbh9DLmiAlJklci4KW2M2NgzgBVQ1rWd
1R2TUmURTXQCtxLUxn/TGFmBZRbks1yF8rcsGR2PK4S0C4z50i9m2MGBUqFzn2g/4Ac+28BVXbcO
fRxs519TiD9slzWRAw4iQluEPWSxliw0JkTzaK1QK1UFS+/jrR0cx4fohnQtd1diaqAGdjfvck7J
wP9I6ANWDRlVlxSqytSg1okrOMdxv6If8+5K8CHmAgTHZDvPNwnnbEi/1KNVJr5vHrdteqtoC/R/
5pCekVkUhdBIyIqeouSQBQHdPZxef/7oKWYuvQ==

`protect key_keyowner = "Xilinx", key_keyname = "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
kEaushxDVdnPYpwXS/FLFB0tvOLAqP8eRXpGS20K/6VvHwDPz73sOGmVoky6V5yynqvT/fAoi/jf
fpZeldqFP5rQtUQDsL86M1fB4uuZviVQ87syOmBSI/5DQDZhhyaE9E/HuK+tX2KXnbyFu+/OVRJX
z0JNxluAk/wCPC+GrvrzBPbf89vNvDKmA2dIZPQhz0oj0LIbNcxhYzgBwPKeHD36/2/BenWRRTvx
IaEfZBrF3yVKP8KyUSGVJLIvxg9rYsKQ02VQh/8L2Dkzm3/LQjcwvzoF8Aj4TwhYiUSmxbOpSBLJ
CG5AGNcLcQPVfvgGJSB2uXgCAmFO/ZIwGKjL0Q==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 565792)
`protect data_block
VZOHbkfRTF1/ZwqzVwvw9qD6eJ2xK7kLS6LYhD1fBEZfiEBgQiMeu4OQUSfRBYQllNLRSco10JuL
zJKqgTuSjTZMVa8Y/mkzD48+Nf3VylO80HN1cEoBYONzUESEiMUujHq3FphsBy1IS7Y9yk3lu+kE
KItlQUXUoKPxpLvv8Qi+YpAAcV0Mooq6qt9xL+T6NihsEjsZHX8537R30A3h0/I+LHyfeUcXm4Q8
dU3PsQIRUMyi9LU0Ckssn3KtngRJUJ5fdi31R6MhtJ8L84g1XNoXwuf+JJiNCpe2urtUO1GvnNHX
64xz9Orh9OcNLOQZnwlzYBHmD4+DUDueh71ZgTCOZW+uSb1IIP+XynOuAwxrGAyx886/JRTmzXm4
RfODW/xl6P+y4J8TNfSct6lVe9BnuxgiOVpLMZbFBEbmoPO/ZjGytJu7QL21AyI6WEtgkXM+taY9
5zITc2yMlHJbgRuw1nvqXXSTjUyLO75xAQ11xhQthfFYiPWURM/fNHv6B36Ez20C3jun5zVHmDMs
jFhzIhM/OBuApF8a4hOHwkgJM1x81p+FQLmDs08Jferch55S7VTqS1nZHbmP4M+0tgHfriPEcXCG
lHLhxiYEYXcG9ZqJ2PiM56ZJNzPqVsQplnKn5c4j3OOZTrznI+mMrddOBSVlmT4ntYcy1VDn2cQi
dv2otU2RZ08LaGHvnMf5uXigjAd7jsuzfKROmR8gfbMHQqwFoIzINftEJ1Pn6iYStZMU6c6jLssz
ShL241xbzLZHHgJ00QdZntxlZS/TNj5gO+iHjsmrw8azTw/3ppex2JnOcE9SM1wnbmnCamuU0nJf
AOyYn1Kofm6bCUqZdCPc0ZYd8q86hzxfok6ByGJhtoBCxlD0UlA84WSt55LkwWki7q9nbu705wv1
fN1uYyr4zaGcNFeGDxRvexJfJrUR4TCzV5K2e7j05DjsS7M27YtP16C3E2VzSdVUVqO2Ao6NbOrg
ZK+25e+of2OLGz0IDhnyIfHtQmOaf/A1+T3DnpHb7t+ZDJVsAvXiYu0X/gytkbHg5qL2u4a4vbnB
SbD49tS9RkYK2bQd5JEeT+tikZ0H1l1YwUYwdGkdkkKv2hMzdIF8f17pvnkklsbtwQiIkPzd44CV
xHWFuzSujVYq1sT11wpvncNyfe0WhAR+/fALfSxSdC+c3Uwuitx3/CxkZxRrKu1lUL9MOTdhi9rG
UvqnX0CXmIm29izftgE51eedOMi+lssSpLNdXq9tE5cF/28sc0P8fsWHwGNZcBUA6NcdkES+4tir
Q5fMXn2gIkSo623RUxVlfoICZ5E0BAeTF8qe20f/5np8payUUpna9KOIU905Vu4UfVNBpMSFzyXN
9WMAPQnBqviuGvA4xYSyAXbB7K8OcK1DIcmpNMNzw2Q7uoVq9pXPt3iXi3KPcQlioNID6eAlfGE1
1LRWa1FjuLhrEQ4JVERGpJrfRlw3dpKpR5wP9DNqQJkkEba26QEoZLWTOKQuSnaYaf7mK6fwsiUj
nk0CL8EHU0HKAbRKwii5O+lCL6plDAhrpaLxygGjEiEsXASGJ8v5Ur5REyIY1WSUjg0aRPN8jK0H
+y0xN9PViYBjCNsYR8LQY+rgk5rsfdnZ48wwJ3jBh5QQ2D9JEvs7TeJ8lURJOhVL8pAVBpQFveqE
KI/2uAjKBuAxgNXsa9WVFHWDrsUr53AtW2gbW7/BtGDjCbDZlUoPli6DO5HXCd2EMSC8wL7yckoj
MdJEulo3UwYnZYcYK3j8vX1nXUgU09w0gcfVwbFqKESJ43rk+MleWKrHHvjKPzTxCVrHw2GUlAUJ
OVJME9FGUa3DaNsNbiKwtgEyPQ49mxnmJjZgJzz0kLMSDC1GssDvBcX02xkhcuswtOa4ZNOuuHgK
Abs6cFqgNtSPeJ6ZjylXn2ev4xsibZmqx1aSRsA4n4/xFrbz55cHb7oc5RjgAz1V82i+u0tnEeFf
NxNIsECkgkPQj54zrG9ucHfPVyWX/4rc9FlQiJIK0mvPq2dgi8wV3TCQEQyHKNC5IHTu7EUyC2DR
xATzXSmtyn3nVGHxWnYW14Xj6hQ9HJpI4DcWJAYzCcKw0YX92L2zCuB9XX/jg1f+pdfxbLeJlrSw
oX+zjpyUQGdWxMYGQA9xUW24vUTPlrKS847c5lil6b7ac2CfiKbC7XR8vsDfFdNlMIyb56J43rYj
pibU49ThUMgnTctn2k8SikAobcoVqE6DiZAkXu7ysXXViHJxajeJqFEjZaISCgCY4zE+X1HYU4Dp
aXzYZJKMrjnviltt7Dbo/JW1ZexPclDMUjd6HEJKvh9KR68BmRuJ3mBySlSDUwMOIRrnWJxFllrK
JSNshHgwEq7UdDCmpRlHgovtrneypE+tkVBXp05Iq8xpyrzEbgkiIjbH96MhCaAoiAASrBGJqZdn
wf2WKRGq/cjh4IleH96Wf86opIKsKq64Zq4kOEdFjhkPCtwLhBFy0oWzbF7/6K8m+lsYJIApERqo
1kcQOe0sSUpGB/DBWbaXjLx6/LyXpbf5VYBb1xBKZg8aFOkwnT2h4wvZiLZ4kLpmUPf1gVVuO10t
1c/WFspK244EA2jTPse4SGCC64UeOHoQtgA+sf4Q6oge3Lpjm4SfbIdFhr/Z8WYrKBMpuleK+ebw
sI30sbkg9DV7QulKETWdJ/yFwqRCzjffsPtJ8HKjrv6hg36Z2VN6cQsBKFlIskojm+FMdkqaeCkt
D99zOQCGEFpCpqX6ATSbf/U4a8BBgscYZsiiOUa24Zlfb0eMR/OdeqIc8+Ahu+rC3UlxQA0iloYs
uWMdi4lsVwucAv0xzkDK611BmkHDX6/K98+KXFnEiVml2CeNJ8OXcyz0BwL1w3wRXf2elFXZ4HMT
XGdStAsPhyP3hmk09t7JvT5AKFi6hml9FnAdWe58guWfgtnWhbqvy4PwAYZXL0yL81AbjRRe6lmh
t2dL6IVGx4JhNfVFT384UuckTvfj5pJ5hmm0HEJ5x3PoTrNXIbNpHBTAGOLfaALvhtfFJFXaoCxV
oJhjdd/cjuqao4sxS4VtYnfeM7MkK/iVz9EmCty2JU5VfSIKkccjHNYAEtqy+/JYzb8j/f+Pti+/
goNCOTUyXcSLr9HZe/rBvHX5+5eIJ2UwtA32OTJZeQ6IbklzC+V3JrmAJp3ul1csUl2+JTTjEzID
zfY3lxaQfYSKUYJhe6UGrlX/R8ltuL4uFsneESeD2r3gOGG6REWMvvs3XkV+eHG1H3Rev4WRdrxd
nBLO7kXcUTRVsyEKi/0me8YVHgcoRknAgyuWROPl0psqza4HKkE+RdKr64Hy0hOuYPUQNk+chxds
970emYAxrlt2UVyuNuTnBiotjfrPi3PgOj1QuisNL77f1DGGoCkTO3LAbucGSPQmmp0NtxPnLUXe
PHaiyylaCBYXKMLli09FQ3w+em7ctOPu+u8mVHxOsTpIczdqI4WtnLQBnUunaCt4BAFVlp4eeHje
Go/yulgmkJAgizoLCa1+tEBPTUtY1JQPDiFleW0baPpgkoDhOKiZd9YoxGmmVze2N9ZiTsKfcxpJ
cz5t2czmNo90ck4/e1vHpDxDy910Hk+/Mop1eZHr3LDD4lnEECctAtoAl68IcLSOilEviYi1GMJ4
85RoH2rZ1tIhGID5tDd5FMMJnY99Aa5/LFV3etxcinZD042dB4iHIRGfYJH3PtZnShrSw3yBx3BS
rY+f2/DurncJHjnT7PZcW5FaBS0Hw8TktwIqvQCApxj6A5qPCyU4cJR0dmeL/jRzivWx/GL2yMnO
rTNscHOkZZr5KzkaiYFysic4SYu2IXwM3qcSFcUgMf2wTpKJiZXBAkXj/Qei/n4W6x9ABWlhUdj5
IZ0dsSgH8gRbl2vcoHmD+uqcBkNJT9Gw41Gs1tWVs5VY9jinf4FsJ9vz3mPaRkJkiVCrYTRQylEz
Ftv1sSXvNworI2QBxXticodto0NqHaFSQebCMAdNyAJPtMOY9M8nlJr1PU3/QP9+ClEsY741fnFD
PXMSOyq1ouY9pDC7Nl8xk7o/rwFPFmfvqcQmVGIUiPYY8j5bGgwU6XYDN3cYwy5MWqj0X1/hQOMy
Gr0/Ke9HP94ExOzOW5Qz5y5k+uRs7/rEaSy4ct0jmUK4h3/SCw1ELatO3BT0r5bJUxPhn8a86meP
3NXD3Rl1vkOTAI/j/RjyMnDUcYP+DLsea8M3cqs7E22G1e8iYBS3VNOb8jDN2R0SOZyGOkk865VF
j4wLhw89wII8MijlrBcyPVDEneMYf+4I+a89/ZelQAGEsFp6nTzJwnkjjYgQtnVWqfGTeNtoD+Ps
hzZ7Lw2leYo7FnRxcPrIOud3NABBzDpg9omyS/kI/ntUDyXnLHHnoPNJDZoVnRzYE98b5b8bEGqY
mDHEfkC6J/U/+JL+lF3XTq2312ak1RVCkjkD/s9pUDd1rAMqVkBSLoCJcIKvOUpOOXuBbBXHhIC9
TcNBxY8el4STvABEHBjPcR3TFepbTpt36i8IhtXu/K7AeVVBWcUuHheMM1X2mjMSlWpYbG01RekB
KAtyokUQpB0BI+R9N1YKoOg9BzS3+fkLpmadfKwRDwQDku6tOQ7rWn2WC4OXsbFrLh3qhSFU5REB
7IO2lRCezBQ06Pr7CFEyKJctApzqXUgJMRTBrdJeAWchHz66GWVFpOmeTsxXlO1Ts4I/yK5WYkYM
I/VCxoA5KB1AMHCIddAKw9a3X4yKebJLYuuMO+MTg8FmDzzRccpCx7VfIwRdBK/IWRYY66GkUKGC
ZkpwJHonR9/YL+peY0USFMemymJmPGY3UOxuBTfo45hbz5ozxyIK4vVBRLqc7XCeH5MZyZ+JiPRz
ZHYUfLeZKkdmjxKRu50zHZqAZwe7CW9NQB1SZH13eEmcD19UxqNw+xSXOju+LpOa1WlZgDy7vr+n
ZSQXtAIVgpzzRSluyA6AtuNKRzN0R8u/tacfkiJPYIFmONaGQzrFKNC3o6NoU45j7ipeaKzADpkW
47OZzkK4UFHeciTTDQBkqdqntho3X+lmEnXwCMBk50OcA/36Gt8vm7sxiXal89FBg9GbOUD5PPhF
zpkW0fg5BcfxlYNSZ+JG33Z73rI66dd9qKvHDHBABPuRxIGRtT/yqocpbDV7aJPbQQ3/Q2tH4x38
bh2lARS6rwBtpyvQAVCbuwpPv98Zt++sVdQmZw/uet3D+9hPpQngUTJXmxvJ9lRgUgF2/7okvHC5
sH5Vx6buEZpWeHlE/IKvfLtT7xUwzp7n5xZZeMA7pLFEVntpGccLf0j1vN6Q/UTa6AJ1T6yW9HER
Zq+KbGW0ObMB42Pkm/M8RzCK5Kwbjvw0FFSwCfvZwphe/d31jC3sKG7/NCzTPRiuPm4DmvxXX1tq
iSLVBrU2vsoyDXADS4MneOvquBXJoM8Ja2VeUcByd6lokUHfwT0WmAJj9sw+uHWRjcmL1+I5UixU
bhsyDMBvBzHEY2lQvtgmBSCjBArG7JIR7LBCeztpDA2zR3sC6ySoNrWA/lf9TV+ryOKaBE03Op4p
LsUAhfGN103UjahPApK7HTierx4IULlEsFNazqQ9qn3re3mR023pUWOxjgvlVvgLDuf59lfcicr5
Z5SfLhQnr4zsM9blmeO7MXCUtHUbC+Z0UPgHS6y+eSQk5oftEQC8x5zQPt8NfFD9UoSH5cUxBFys
Atkbx7NBTpyaXMeXkf7ya6+VT+zWMXgwxnJJRazD7NHGosOJY9YbC0k6RJa++7Sm/rVQgDiXlmxF
RGKMq2/1BEa4WaVz4OqCRXxbLejA5PIQs6c1yPEjng5LAOBL9UdpMIUrumd8Qg4cqliTJchF3du7
nlOfpfZVEjIBsXyQ3lkENFHzfpwqVqmdwlWqOLtsLfUbMkdmWOlYy+i6DPJsYrtT4xiBmZmln8S2
rhVuHCLAiJmQ4zTOvrgpO13R7UXCF1m5rDldb20QSvRLWsW8jav6HiwxgoOGwzlxrzXCi9L+rU2O
8Z1y27p76xr6EzETPmNtxJ/+gr+3cIVhWl80TwjDCcmD8ijL1tREFcwFlqvn52LILjCDtIzbiSSz
3f1Q9SADFULdhbId++zCezH41CPVThSUNJFtUlwZK6UUx95w1m/qAzOOtWEMMPNb6hHdlIrxBZWX
gCgo3thnOoTSDxYI7HqMqY7jR/x27i+5/RGRaj6sSlNpzfE1bTOLGUOwiqDO7fxJanMsKx4fOuEq
Ct974qAstYMzy3z1wMKdBoYC6YBJDPF3DbwQuYS1okwwsQZvW/Moeo5oByKBuZJaVHTjiQtZdJiH
LuzbwaF2KL02TLWKZfJY7TK5IifM1IdCMjggTUacNSw+agwRkT5RmQL9gJSnjCLfGl9oYQu3zBCH
uciOlqAJOuUFLu5ZVXwUu6iLrfZeQKna55qQBZyc3BOIWiiyA+GHCXOCoBm7AiWRHH4O9OKWEWmo
B5iVUn6N3P5uDXz7YL6HnBOEYd7pUfnp0/utKmDC6Ba8bcexJMm2+yMQwyN9rxI+sxP1yWij4GWf
+UsvzYuTO5To/7pz5wjb7JFZO8Y6+vRc0YdMiAVctaE9uwFJpnFM2fquMQr4RnY95FskYtGmYo84
gGCuIzadc2MQQgo7nW0mWkqX8ne5K3cOWkYtqzgfvjYN5XIP+Lv4U8gMkM/AN3iV/u8htEXuqbhb
Ro427MHHEM+uJ4BpzY8sx837SuXBVeu1scJRwuR1/I91vdXFWbV4iZHmS0AJ0342+//3RgLCXA+n
dYquDLHDSGL3KNfQLwazwsyULWC0ONku0jf0VfLKAp0ikdfteSTqdjnyAKqCZvyeYw33YWZqLwbi
Dm3MCAo1qftJB5n7PeAgvNe9/hlJduJl5hxk5wBQdTWwg5mmuhubym0LlUjBC0lksrI3k9qX+H/1
x1f7fZCAE7FAJxVq40g7UsZ4o915q5WkuGAMBFVOowQNmLnBmeNrAPY+MK0Rtv42qZwoWmQuh24I
aKU7dVvVMUsEiEIJfR54KeMgZJ1QiCWw6UXPfTnN4QWTEqcXDDJt4FUCvTjuhrUNo3D4fuyyP6Lk
TUwg3FMjznXiQIiS8yzVxu5g+S+6zN2vP6v6ffMf+6TSNwpdmFEVu9Wh49bD6qIYLO1Y+TW9WXEC
fFPTBeOeYZ3iWD18YoQHRpDjM6zWLRhb6cb9SsAY0rvLjqZ8l2oBUb3lw9jgPa4NzD+IijQBSRLm
R24iA+3Zx/L1KjVPdkpeZc/fgch6vEjkARIWc3S9TSmQ598VThunUJF1xyYD9+cGg0qsV2GVhf8E
cUY+DrK0NrHGZCMQ6Z4/euL9yHKE0IC44FL51jwDrwquxp5p2clDpOYDf3+hUGhV1SFuDpQ4VeJo
/8R386N52Y0PfaA526JXeRDW+pujy4HndGzpwO3Bi9iNS8ktptQ5sOTXaG/1y9AgnhM08r++sfDY
FX7p5mlqX3DagAr+xngAJdwZm7rSiVg8z89yULlkfP39FaD3/BQtHjem+vmPz0xdkgKffAGm2E5s
x36ufkeI3o5DRJDrimds2hUrbAWgZw0N2TPpmFW4wQXbv5pl3MtLziWQgFHhEqq8f+B/2E5ykP+7
AUuaOszs8oNzkchSyXAYfrdvdcSqpWbjKQ7f5jyoN4kLxPKcXJyeUKXlD8Ji1d9B76n8YqDmSk/d
U1nuKubxQTPaFBVRhLtZzKrZypy2d36N4siHBkgvef+zVIuTWI1Z17ab+hmIYdWdfzywobYWg2Ld
ZehKmY1fqoxbds8ejtkTtU6kY7TP5+QY0ebaufHi4BVpdhgnE5xt2G/Ta9kHXAeI6bLUJ+XRNH7B
yPKy4NmWiKWcHaU96uyOR5eIMMYwZ/bXjytTglVCZtSQYp8bmx50OIGlqES9G+06OCoUbuGHaS5D
Wpg+Q5Zn20UYYxJNOfATADVbyhnWzYs1sIAb6beg3k49/88YVrnAU7zjvCsi73PgEn7sMuB0dfnh
/nEHjccQAJjyIJuqIgy1JzeshovTKxCAFX6ScmOedyi1JoPRatfA4D/tlV090KjUVk8g/GRBR4/W
6rvsooRbeYTf/rpq+JY4Wl0lAPEU7ONbfen7kIKLdFOrR+pj38ffSM/bP+HR7HhHi0ZwBMJolbCX
6fZ3YPEjcLmTm8qZwcouaR+KNXtxCsoenPN62MVMZ/a5sIN5txMC68rHJgOCz32xuqJWpsgu38V9
eRxOuw2X3NvPWk8tULnNrI4Hqcg3E9nkVRDp6VeMTI3w45e7eJUQPe4Mo2MNYUwYGRjb1iUIQMxM
mK1V7b0Y0+JPLlOJFev+kaVQ5p0c4JNB3jYtGZ0KditgE8HmsksIKCSGGahMtKEoXJlSsf1j0uEI
ldbTQ1lj3C9km2fAJcN1n3tP5bFvrb21kCpQc0L9f0PcYACy90rGAWfiT0ud4CMtjRPYtC7vYD03
gdyfRu+ZS6MXvWAIj/7lDyE1UOz/olS+BuD/L1sgNCQvg2vzlmsZoKzeEmKNnZfNVSQhxsNEVc6O
d8y/V8nCEMGZFu094NAo6+APj/FHcMLsqp55qcXuTJfi4DQJsBLIjytrfXlcJJbLRLgpYvA5iS+9
2usL4PsyJrV/breDdsw6tunCBIIgP+K8qmgWmIiPmar2vCYTmQQrCl/FrSyXkxbDEgSUA2iFJq4F
E5Jb5cUDTcwvRTiU8ti2SUl0qXYq5a+EL9ri4nqZ15cpcGM97DRIB5ZyC888c4ey51X6WrC7yf0v
aECvZjLjKHH8CMH2Pm0zx8lsfh2VVPZXJsJ6P6LmmHVVcNzTvRNKz28pC7rCF2kHtovkVqVplice
4nPErRGc4T2Wk7iofphbrG+joF7hoBSAod5GL64hFSdJy3/PdJ5KjyKifokE/EWEcLR3xrGGWdWI
oGFgeTDXnJPV0Uz4nhYEAqPJc/QOlns8j/cBDH/n8qq69IoInustw+Ej9gNSKT/WexS7BeZOixF7
UcmII8TQ8iiuqJ3NTsGzAd26MgdkqsPqH9sH38VQT0ogNSbCiH1QclCQnbrC+2msd/SSC3EAcy3L
SyC3eDP1fZtr7HAjQoFSQB6x3NvdZtpw7P88oTgXVA6IZIu5yaI4pS+Kb/bqPPosQkJ5FExLUHzG
kMsrcroGtUrZzIKgeenj/ThIbd0A+fZ0Qzz+VxLjBxsHzMwi8Q9VBeeV/NUzS97UDch4NvlmNcob
4R+1S2xeG8OuUWiZIK/sxU47ZpKj/KcQXIfzGreOknBLXxPpd6acNwATalX92MeXvnc0M0qVykh8
f9lzDZc6i5u73hxz3V1G5OPew+U/foFglLTXrVap7b7P45snTkJZZJg23B6nKXl2E5A4ZpIbYP0u
Z6BVObikr7KZddpr3vI1+lRWyKSti1w0BvaJPDmpdZUvOV3ZBu306xg2+ZtsRQui9X9EcddtA1Gs
4+u5dqcmNTvgVPSKie4B8AxL8MUf9FBhupmcu+e6NE9Y8GCpGs6djqAHmW6ZV49Oz42zFa8claz3
BhdaUt5QDDoLdV5er6tRxKq6kqdmh+8ZSAz5x7B5o18rXZ5ce97G9aIHezvTn+DS9ES4BLrGch1r
dII3m14UV2rMOKohdM1spAnmWqOl8AEX72e+vqpmPOYo+JQmFAfpxhl/eROdIS6U9bDz1CyOIjG3
p1KEL1I1moSg1PG13/xb00rOQsJaasa6y9Tcd7pBJkUxjfiy2GU+Mb8BvU0r/F5I0MiJnx+mVYFO
q1OhiqWKYVPet72hTEtHrX4ToeBU2OoH2XMhNaMdQs3Phl40tAWqNjygHdbN9P1ssVFhDFacPYVG
pr94Zczsbpa9AVlB1S2epOxfKzjYjbgkn1cqOrtpYScLBIoDeL3R+wh+LHB14nd6LOGifSUMznF8
rMR/ZiXuisn10oY9n0fmgvk6tTZP8Guv3pOs60pmhh8UbI0VMGlCE5dxHFRRHcW0FIGqvzApbFM7
xx4JAIKcN1aQ7V5R+bV4iNc9C08BoL70dDmqIVfbvBI13U+jgaieJFHWYrdS0zUMwSROJ+b9hVf7
zXB9J3pDKSjBiar/sj5MyxyBIy2sFDX9WjLdk10kxF4u8CWL2BCsmBnTBv0w0Cjsv8cfJ4NZAgLV
B8HnV+h2eyTGA18KwD7bz++OUHJ5Qs2F5Np23LvJWSo8VsAmIxO031TNYaRfcK3lTV7n1CUnzUfy
uSqWdTfvUY18FD5MCcXwjnDN5SJ5FPWHRRGMKw9dopnvSTrqsU1URj5grYyQxO6tnpXIA9tyoLup
riRWK/g26reCsveLIXZ4iDPQqRqJvv4SPUIV3hXswSv8ojlMbTDs3lunSeKILlgKxbPGMchVekVV
f94qGiQUGClR1G4A1MMgI+jeQr2EBSLaHvICWgJB25Mb3fZEe5YX7KQ7c7Eqc3xwumYDSpHS8gdq
gE3wAeUWyY2eOjLOAU5NbJOpUZgog4QPNejD3Sr+RXLctxjSBOJG+Yg21aYUiLcgllu/9WmBwyM5
woXcpVHkDWl8rMlhhkHhU5hXEyvBdS3uSkb5j74r614a09cvLFhCBCaVR3AW/TdS/ZA9jgonTuHG
ILDZo9b8qmMGvLoyMRAuw2y7hVqHbXi9/HqzQZL4XPreoJwSh2tHsCi/aXwkpSjildvwGfnmiXAX
FH14MtQeZjznOnPjMzm97yCwLqJ93LH2fwuAbp1GVxsnZnN678T0BtP7lapUCiEvE+IWtSxliZsQ
IpQ4GBVTb/mqANYup0qU1HQHhRB8MBoAJB64J9iNSGyzztCdn64uHY+m/y0LTrK67umfJszLWkeR
ikt5LieOWc/i7WdUXkJz9TG0g68PqRqiN4jVuoL+w66b0wGrfgvDo6wsk6ubnSJf0qb9LrhSvGre
jd344gkygJnj1g+JYlYR7XuDNBfsnW93Pt/bpsKABhhHd93fl7ppLOxs8if4tQl7e/leIOYM3D2C
ePcBuY9oMzO7s3rssAWlL9hd02Uh7oOUFkh08wUGcUjuiTKCSFrxZyHwnbo1yrwNlGjTjl/NYpc5
sJQ7UN+qo0czOLeN+f6AxiQXVs6TpIQ5HfTv/ADTNbfQ95UAsxRYlk91PzQc3QKFtTG90MJtf0WQ
m/2JtKIgyrRhBKbf4mV5RF/m4VY+apqVKVc4XKi9RrOchuSbkaFH7n7wHJGgM3DSKGjUMw2GHv9a
A/S6cT2EJehcFk0Wbsz7K7ecAG0WT/LZr+xlFqBuPBGfkGZblQKC8uPK1/gZ2zFRYFbSnKPDH4cE
bOtOTdS/AL0mdwRNUTshuAEyC8OacQyiBT7Kr8KO8ic2iZnrDwWL4nIy+SNN6EjJYGQu2vL9Jzgw
H/Rn82z3WQzEUZLnf22NY1T4oFgAkVZYoMAES4v15pLdV2TD6RUbH8FEJGe/wsJZiJ9zSBjSjarm
sJHlRfD6KpEGorQzKnQO5tTgH1uJXXQdGYcrLCqJm1X8IlLMmjUAxGgW57JK9zOAnMQ2fcANAkfn
jcHzmHGbqqhfDCskE2z8ANmgEYeCCVBYid1jfvkpZr7j2I+CTqPhX9vW/5rImEzk41MdgUHIroSQ
caTr4Kb12TIJg1P7iWrQt+9Gu4uFNp4VfM37f69uSAN+SCgaeajnTE9k1ownYsGMSxWqtJzz1/wS
iS7GTL6w4z6JyFSusCxUPkesiX1tyo76S1b5PBZEsB/gXI+e98kVwOxMQlPFtRxO3w1snohhLT5+
T3u8EoJEJye6CC0/pZBqErZoqnOKta5zj4W1mMbIKh5IgdOnIjDdSs5aBjDgul8FyBzkX/x8eYRy
8a9RuvdsLFDtfoA00GB9HHSbJ7BEgbLI/aHEPQ4eqYdRnZB830punf8Sb0uppg05Ldvap9L2A0FT
2+lNfqc4B1+1wcDrV7Yb8fpp0pdZGfad9iG4LFlVBGCXbKMQAU1dDaXUWu8ZkC//V0litrfMiHC+
6ZeVnA+XHy/tvMnJ7AFsYUbHaFXM1wxQjSfd/3iTsl1CtiR6uvq/sq8uvw7wZbr8mpIiyyGH9d0K
wqK9WOMjlDKCEX91f4Yef2ZVdY/6UH+prE1aY1rvwX5CZksxqndof3jgeoJLnw23pLsWeSt15Bcv
1l9aG4iM3XOkpZQ8BJEouKh6kBYTDmieAiIq6gk8DBe8SpGbrSxAS1GJWfJYVZNWWo7iFlwB3Ego
DwGyMbjeHZQGujPgHyiTQ3vSyXGlbbr4DDH/0e0lYz4CnvSu4Q0ri0s3hm2R+/6s/xJIG6h7T6Hv
Mm+rIsSKJzA4h0J9G6GhebUbdRrQI3c1Nvvl4ep93kT1Mb2Wk34fTeSayfiwp+XOU74KSXJE29Pm
YEYSmfNTzKIrF6YJ5wv+XjWUN+WG1ANtcxCGLiYPSPR6WwZBxx5TUA1tjVttJQ3pSWYbj0gMeFfQ
h8SNFJYsF0cI81GTJYSRQoa0l9sP1siD4aZ1Ay0umSk5UTWeCpH0gYkhk/mnmYesEkcVUyVmWDV3
kekKGfnvozo6N/MnVIkqV//pnrLXgtB5MjNshgqPXgJPdtOB/prDoEjmrFkqHEOsgV+iYZgdEY8p
kNjZUenJubZXjlL3ek8nrS7tV/VDpp6ouqehlIUaOYKcmCUMwcPHInNG5b9HlGtkwoznLPavzfhi
ALw+/21ihq3gNy2D+ZmCvaB8Qv/7sxP8IkzFYP3p2qwqg+xmVBXgUElJShiDNILxNojnTPElfyjt
bcBY1RfIBtsfEiHjPHCO8lmnf/xXZFCjQwvHQ8pvFpDNF01V9waonVJWZhvoY1RN7Yx1oOtqXSyp
fHQoaR1egxOfyXLM8ABdz21q/Rmtu3SlIGVewTGpOd2aIqickrH9u+zwXbTh39bU99JPrFgJO4Y/
j8VFefdKux5OSz9UeR7ok1ot7+P5pkjeBz7jsFtT3qi4fc4Jk4clPyCYZEWNf9PDQnjT7tbMKDhu
MWMAaUS9UdOwtDoNB12VsJ9mcVdzC1G1z1IkGObrGjY92LibVNm9KcHfoMAbRLNkYmrj6NDkOAWz
wp0liKhfHDheruyijKwoMMZji5lcOBEmImQ3bQFuv4EVVJcYjIggra42hZifdWIuGdQJb8Tmx2Mi
oSEPHM41qgSgQMS1k7MrOaZ722W2yqOMN0OqN3okL3cF7MmFevP71lJEz2ERYwKOaOxZ0QTYJVKQ
zOEJks3Ik/t0yzAZgFYghgHlg0XQNdMSAFfH4kehMWqEtwoU5j6DqCfhFUGWBAfcP1+LdGPleMVu
Ne3EwvywdAxOoYkvN/1BglCUnyLzS/QyVGA5P94wMY86Ctl897CpEkUYMsrQPd+snFyINNlsPIej
O5cLJVz4imO0S3G4z8ilIFqC2i8JKXAUNniQDaJgUw0PE0O3tRL0arxheY3n5IVgHliniLXBCR4b
PpY1cuxVZHNInjlwq2/k7+voUGnPzPTHB0YUottSqmL90mM77Z9t5Fqcpi2YHdmxiAM+49cwB5Ad
MqZimWL49Z0vtPieNUMDITQe6q0A8p3w8Qad1iIGOJ+KhPu4N4vDfHBL1UQMoTxDuxdumZcvyifk
4oX5gDBXV0rLvIdxCgVDzJMgVCY3eZGKK9Vc8JUM4IECZIBb4PWtGocbDul1bgnDTpMKh/ujgRFw
KVo6SXedxLVANnI51/CjVn9w+yVs94eGKHDjz8wKkCrXOTMb9TXNsfIaJRvSVavAD6FubN/tqF+Y
hRSYDFLoNE2ZSbCdwyoDqERbmP9HJX0uVgNoXNlW5M/IEg5RjZHbCbe0qQL65LkXIFmUsPtBFnS+
wrTd93bC6+jmsPdnRbl1tl6I+B31JHkaawQlGyhkoQsbQ93djwFCjUdFW2qC2qRN6ziy5QmsdhDb
2jhFd0MZ137/EEquf5wx1B7qTbLP8uTPG8TaIqoRooV5ihCjci0pbbjmS0TJdW1gsn19nfPrOMyo
lSW3lTfadkXjbk7BDIg5qxk+/mW4iMyod+oVhCntOMFFpQt0g9FNpB2oP78NWpW3K+EdC0CcUehL
KZpNxVrx6Svqa1PlvTvoSMqmbMHpRTXd3MOuOT3wZBm/VFj+J8qbKlAYOsGVO7tJlBG67hV8zn+M
styCXN6CDQeH9Q/qld0Q9QypoDaj918VEsMpzBMaYFSYssKWTyZLeb1/0mxmJgc6D5BjrvKV305D
67my+7DAahKTh8gnS9XGiKImo45hcROpA20ksqtoxouhlkChRdZv9QS3XGiHoBRudoM1dLGy5Xfd
vDj1+8puE5MDctlUdT9h9D96IIXzJUDYLwy6cb3DhV0Ula7uyk8ScmKxd70EXi+BOBjndBvaxBat
C5rIKUVpcslTPuEoznltWIvbVL5c3GzT7DOTHUqyxDif+cbC2vccXrdt8HPoU6WscEQvsqSKHylV
1b2gXQhrKxEDUNa6EvrrDmacIzEY0ChnoE0d3go89AHBkDNwrQSab6mtjIy7uhOhp2BHPx36rE9m
bUPCRFU/y1uge3iIwMDMIwwb6f7bS2EckydVLI0gIP0NTH695OmFZtHYC72wMRhHDUT+nJoqdHGa
odTbm4HcQ/Dw3mTzl+HqLrHalzB21Ef8xlMECqsNK6t/zUp1N+QdkxBqE1sIUS3LLYaU1spqV13n
IhVAZxn/7oGaLCu8qVTZ2MA4smi73bWAaC+siVn6VbB8XtJUut91mf6RALLE2XjVziBOJRGdrZsy
AMgPtqazJwfSCNPMYSa7y7g9ABQnlrc6h3EgcVZMHw1nqIJlHT/o9wUGEpxksYgd2jQjhwCj2m3W
XAD3kkbGScvA/kaxRo8kin/Mlq3x4uyQwkLD35d3VTVjfGNcQuIzALCsCuZ7Secv9oEDEm8yPXod
/Vmet0rTJj3GzLrIhNTfXyaUsPtAmXRElptffseKMVI10NpXlauoNaG6F5QTguUnQydYmB8gAyTO
+meNhpeWrvPt1TY87+wRvh0VgbuI7u0ArdffC/2aBLazB5Agv1j7IJ/skfNvuSdbhMFk1Q7yw6Br
0EoHruLT7+HDPMoZAQRi7d9+uGOCP5KJayQGtXzrll50sFnQTef+dEQq7Nhy6SFET74ZQbirLe/Z
YVlQV8ayDgkAh3EAfsnuaCgucRKJ9/5H2oCMks6OFgGXWojhqhYubNGDFs97xayk7KmXxPy9FPKe
jsxr+1p0x7gadNOG/NsBwxQEgcJEg3/Ds4ikAO7wS/U0HLDSBol+9Dcwf3j/x9Jqe/UPV33Mxb42
TSq9Im576ac61cXeDZf9niaMaTREngjTN9W7BHELQs+SJ349emCyoktTq68lHpgBndm4IuV4jl0W
j3SqSS6n821eTWagxlu3GuffRMaYn8GXyykIzsggZTF5EneYQLPugvWEBd2PqP4g+6cWu0Ymug9h
kIv3F+tdmjIj9AhnuiwPhQXbZHFvEdNaptRwkt1woZdDZjqu0Ic8IRxybriAk2SPW3rHMakH8rRK
vs7WDHb3VlDjoxPoQDJST0uiNcnMpPpbWR6T64D+xlRgu7HJohCCK25Fkb+BzANpGRKjx7AzyEMK
sMIKajgIg+SipTFGI8nOfqzPdFRr9/mRetXQb3u/nWZpprZp16gqtygQlD+5d0nPm69SY2MUFSXX
Q+D36HRobXmn4x5N1GBxGUN/BP5ydbWWRJltZx1hU46yeysFltnMfKbF0x0k6BGtIwt+rn/wKZy2
6QhYRtZ4qBT6sO8D/d6Tiyh/VCeMPbFHTcERMh8/BW+Uh35qbmdKhSjNEY79yjZeJwhBok5l+Qlf
1Fz5sX7MrV3p1y7UY2CXlzPSaEp1E2D8ez3rIQ8+h6cnd2cAxLdLQRbxgINb5nUuF/aB5lhZv3JW
SP+D9dmBUCibRK3JPL+sxUBWeiCKkUw9HXrH/4ea/MHct/IZIcWynY8HaB2s5v0G/O8G4dxTAfhu
bNw3R5QguYT2Igut1nAB7tDEk4FbvJA6fCi2TbEnyMNJ01Amr29ppOalXlPaXW3+upOpV508UT6H
wENy19F8mVdUQflAdEWDSaB5SU/WnXq3wKjLkUT6mpICEp0D1QB/I8Qbs1s5i/tl5RH178VOdLuI
A39uWg0+Gb7GuuP6e3O00Q8NBD+q+iHlUJH8tFM2ychVSfk821lZSL8JnVgwGMev9rzCuW3JylwN
VYXo3QzCr8e0uoKTnwPynMfZYViql5rd/Ox4WBwVIjJymtjz0yMpcstvYi9D9PgwuSf5BxMHkcyj
dYofwV1KfEYsdfpr8orYPN1CmN9efmrGJxIaiQID0kWOCefy/KyHpcjDGzatjYZmjsPO9lyXc0aE
t8/8owyHZfiRK7YBPDaK7Ga9MwOYTrj9sZ3bTwHXy4MRtiDrFQqOoHoJhmi6YqU4HFUaZRT5LJks
oogA5G2AOmiLrYr0q8KyujCZVJfZflte8lOqZzJtbhLVt1t2wsn7sSyks4OUXBnq7BsT1gNxwPGe
+6r5+84FiSiTh209Z85P7yDrkmDnbWSkpREGUurZHz8Nj7DcqNO1PETp7LMe0SWS3Aa9sNVqHw04
tYcAAwbfiCaFLpxsX4+m9J6eCJCOncokL1Wa/0mJY0khGrcIrd2XRPAoiPN+VZydNwpjj+MkQoXr
uB7UlNl3OizsmI1wM3oIoXDR6qUbVLptZ4m+2BVW7BiyaqW5wQMG1WkAkGcaoSuCvN/39CwQIUGa
ykICE22L9kNmdsAzGCxtGyhCNzDiAEoJD3FnNm4dwqi/SsXzL5EIiRNVKTRhrP9eACFkDxJSUL0j
4Qo1uki/XlgV1QU1D3THtADCiBZVmyb7Vhvl3m1/tIKvXTG6VKIbeRJvTNQNjPNFHYnds0hSFfnr
kITmIL/CT2ctmURKtVXBglKbCeYvxjYx6WOnnJqOZN3t7OR36U7ZntHv87SZJsLIzY53UUPAn0Jw
5Vs4qNhVkHIYkotgLtU77za9Q4FV3STu+zJkCrIkgBZBcOhJs1lLpIa1Afek77SsYIY5fq03B/Ms
ZGvxmHksI+sNrebVztMcqAW0ug7tldnNzOjUHhBnqHWB6IqZpbvplCHVkR8ud26IQCbFulovUDqr
sZDrTHKR4YvyGPUimjtlwOotUiX3BaB87i4rn16q14zZKjVI3PHjXH2dWIjYDgj6ni6UsdGw7NKc
0Cn8wcXF5wAvmLCkF9BY8BOrkqXussP7zf61xBOFVoK488tkCL2mQXI0mzMymaTcbyQAIm2hYgIJ
TNEdLKJdT0CogDTdeHGMP9R+KS9SUpHZkExo8ZQgTCiUMV+C/iRr6De6ib8FBuV3wFaLjntyGHQZ
hLIzloBvKUL4dM0hH8yxyvi1alBJnnxqrm/SyYJ7Py+eea4vs8AbKj9AD7kXTEbIfNLgRZ7XyK9E
sLFnjeIleL4EgFfmaSUgpgWkLXyDjoStifrwyCGOVOf4q6Wkfec5mL28DdH+1lJFrCZ1ywzfRkQh
3R6eMIRKzZZfd7zWrED+E1/v559+RXS3Sv1Ez2WvWju7dYkfFCzJM7STORFsdChv7ZfPR4OBixKG
yUid7olGSUeSNNgP7KBPGMgRHx7j3OYTwj9Dq9yCQ4UudHO9o9ny5WXuUZ4lGNkC4rGvqpJpzVuB
ZmOXLjFY5UFMcRYT3xCvievgBRnttp9lwEKIKrrRhqxXaEn0IfOym6t6II+mrJhga6z32yOl6Rp4
wYcgo1hgRzUyBJebTcgGSm6ezGESCSxYHMbwj51WtzvyUDuBO4yWkAOuJdVGlVpful+SOcRnql0z
YcDbWKq1vzjo3hui8i9wpRXXhtgGBvaN+tccWyRfELHYrLn2b5dZ2WmQ5gZoz3/7yBABG7Bvewfo
OqxWdLhhfFuys8uEa5DD/XUiapYn23CE18s4UGuZWm75ON/pLNGGVQh2DGSkRyOi0fe1NqeyIi+2
bH/+2YzCiCGzUz0YS69N3EPsYwuF99JIAtmmlE/qYcu9nxn4YXFvWzPOWWpJJZvWFtLkwddRcDk0
/inmx8K5rqpAw+u+SyyyrFVI2jBYD0FWPJc9Cui8bIPP1MMkYXLyTNINZ18UYHbkrIF4vfCbdU5o
pa5gNKT3xgqH8wrJUIU7Z7IGotZzKKgTwSTH0R1Nz70YVhSoKbuQ9X5sQopFVzTH8wnDCTpFzpwb
UDVFMWKXT2eHX8iAN/gkRW4tAyp82j3DBKkw5oi2DQem37KYJlCOFOBtGSdU25j08Q/ZH5P2O4OS
3I5MhaMqvlHc3knHWQBc4d6l9xGeoc5GJwEVA0RXpeB7Zeb9xwZjf4StrPhdLDOQAx2T24OJX420
dN7LwdAkstz0ZCTPgx0uY3sq7GexnjHyomj/6Ro4dSRUFT0MF3CRU9xvf4a7cmCUGtpROsqoiw1D
TcTxRlfVH3VQjZ3zoBI1XWWq9pBbAaUfPyV5ZRjLezJFFCBjomZF+vwaTvTqBt/gFtPnHH2pLewo
d2UA97WVZ6OsSFjcbtqPm7gCBRrPiOeNgxe35YMpfZVSIKySiaS6TtlOrcxR+kEYJ2d9TW8ZD65n
q2TF8DN6JF9so1oLVou1bi2LJl4lSA1J44C7VWBJVp0esawfZwDau+u+0RpGw00EtnWYPtnW0hzD
0S2f646K2QpvK+pzXiK4oNb1oDHqPp6bvY+UfZ9KMpGChNAXUyMqniaJwRZbHisW8iIzCUK/fWNC
u0R4vS2SRYfU/axKet8N55YgKBmS3nVMz55Fq1eMlWQUvQLzmzuwZlFQ6iXdyjZZMhaj0a2B5bL7
ducfDovJf9+cz6jRB0UfRijOrGHCx2Ts1FyziOlVDGU5gAW7C7RiNo6DrIWc20Z0Mvz3ftnoq2yW
i95Jo/hx9foHdqBwau6mrvtyrQ3vLndPo9ZbNaMKy9gIm3Y9ePBo6F9ZI64UL5gxIa1PnclgIn75
jniG0pxXjkq9ktx9eQ5hCfiqb7uZQDaIzuKom3K5bheuwsp83xolOc69jKbyWsbYXt1EvAunlCnq
bNSEss3sr2VNv0KwSV//1T61v7atW0n+2dgELId1bfuyrIKj5bHU9m3JtoveINuf59xCycPJk1qm
YzZ232Va5u2nFjJcEZfcBtU0BoZZF23ermnG6Z0HzI6KXFVJWWiKfDW1R2+mc+Mvp2uoj99eefJ8
fAJd8B2U5trxL8Ax7X60O0jNYGWVZkduajjjMRZGGaNdxXcTSY7X6ZLpU/xWdkJgUViuiQE7KOEU
d8WcVVy63r/9XEahlfxkume4i9g9eyDiNexhc8Xjok264mgtT6sb0zNawpubmQoI2nsxE345ehDw
OU9uEe8CQorpC2wvdefIIoSVcQiRoyN5yohBU4EORkr6fLEJopCksCGuAT2sOZr56htenMaCFIfe
1jj/STUmp6FfeQeXcMATfgPR2fcdRDY2GDb8kP/PtXUU4zqM5cPueYuPQgB6/PzeIOyJo6N3iTlg
9Ga9fTXPEZQelJ0uWIJHEv0dRLdOI50mxmMxJSOWkRoD15i2Nt+p2MUxoZSpUvoeTW+EqbRvjIUK
xIOnBxqRHgVQlVATr+0dCqINA3mgjlcR18IHLugMOxOpdR/KDhwQMgisB8F6tAGcPnw4Ats7jkzM
dc0zJEdsl9Ku5QX71tjtfHBe3hBFH2DCLULe2BIYu1bTZEP3gJ1qdypEa5A4TdUHUixzH2ierH7l
YbufXdW1ZI4o2sMFneQcew4ujt+CdgTrurpuyKVCMQn/R3ORDmKCTrNm4xeYD+UezF2GeVVIJsF5
o6QheYrkdOvnlW5A19CU1Xl+YFpyUClaZ9uccyvZ68CWwiThssJ7dtshas4AhlVARUE66+sgXgdq
xZBp8feMX92seS6UnCWWi6xRRAONPTBiUaNsoQVfrN8Cl9LAhmuIqRQJ265Kmab4VwXgbrm9ji/f
UwUrE1iBOqXEw0azF0pDxDxqcTbgE0zXAVkAnpNUUxBJympWzaeM7Cho1xsCtrssWYsFLUnuY1ZL
8z2yMnYWcuCRSv61maeP2+NodaEFSODCGEVMX84aExj8kq4FT15w9KE0KDZ9qAA8GFxQYfiYwZ4B
5yWnFyOIOBGktfeUq2Y5zKhOl65YGXyEH5wwzgxmYiFhgIZjw4EARqVSjL1THVigP/jcFkZDM8aX
feMPyJueS2Po/EGHhPq44wz356KIHQQzC+oveH7mhN7IVdQZ2WSzn4Fglvkk6IMsXf1hg5K7HvK+
11B6Oj0g/uUNFCzte+8D7MTfFuG6SMlwefrSGjiEsqiesIPtnb2I5KpLKVuWcB2hn0rru6Fx8f99
HSYYVAEUJizBP8+uZR0PLP12PgnxIFNDNEaoN76vu2c1CZ9HQVFojDMcI23mnIfoSY2PnE9QgzCk
XXXQN/4V94p2Olm7sAZwpaZjrjEQgPfbuWa7y7jn4zMyIT/8WIOqYQj/SKDj8jGZZM4M/eEVWa3j
jbs0N8MWURzyRKMYrl7EJsJF7z/7QINulzF18qoUWVTp0gBbVgwqiqCGXuGQ+0nEYD6Scevm/xX8
Tt0ISemAlnQ/2ezXPF4sNUkGaVv+WpfN9UWgustHv3cGU/rbYzVGItsvntp9+yJOM8LUjWrRy4AY
tUJQM/5f3USXLgg2gBeB+AoMNLFHm3KugNfQb484r6A6tWzerDtS9qUnec9U0Ckr4J0TqHRRRRj7
ILEaX3JtsTi6enNkZ8vvXWcWBNhSCY4vxVYBoqedclk+NxNPiBum2qQWIiRpbGEL0tzCWBq761wk
CI0FD8LRt9pmrIm+kCr/EO6//Lqpm5X0P07dVzOGRBZYDtYunQ/23fD6Tk2hL7mAIncO43fpUKte
0ns2fR0eUX92f2cL8zPDzj0NV/CLO8vss6SbsObKT/713Z1W395bRpvipVeRWdxhtZo0yKPrk6vY
uBOljdZxO4QreBLAnCiRBuaJj55NQYMDY18SRP52h1Wdx62b8rB16PAvp1o9Wo1knTDCIw7MsN1K
jx7IAvGi2ksFbGMvAE5FNBISUegp2tZc3a1I0EmkfjC9NrU9xZePi/E25dnAEHVZsx8fgSnVxcRo
Ui90aAIkWoU/BsoauI33ZqxqKwdlgeMtnRL+z5nVQD3kwl3B/unIDRFKssG2/9OPkOYzmh8E/Evm
O2v+QRawchumxUfme80+ovBTnnLZ4md6SzLvdb838O52JZDX+qL5D4CiPQqY4frABGFDgAUnk+fH
WksFAUOQIJulvr3zPKAYmI09IKQIH7EOPnEdw81EL5CHPuY424vUOSDvBaauZOqF+dMPMN2B8vpc
4DcJt/wH7b2mkmQ2AUJwR1RVkj7kvQvAUkILLjcu8Cu6HwMyedVEAvU4vSVyh5xA3UrF07B8wWMo
dvc5hM25FyvwmHJySAGDmnhPNZoeIC+G+El6LLKcnD4RaA5yzUjonsi2nzToNMwZEkwm7gxJjzAW
UbeJyexG09zs3m4/nD8kkBetfl8NFhHRIDaKCulI/YDMayRGXnmkEA1OcnIH00PcJAjon8Usp4BY
DHcoAdhquJ0L4/yhrVCUxQx2HfkWJBqvUYd2zlpIoWW8G2pf+pdFXhxMY/fIhqNVxVwr6yDX05yr
+CxJ1JxNzvvAlZukk2NGfTY14WcQNB0kdpAIwaJrDdbrNowkG4X6EmDIwfIEYtJoP3y4aJJ1enud
ZCS//07QEj4Lzz9BG/jYerRPysRoyjQA9TN/0x+KjMGW4mO7poI/MUZEU2dS9XqWODmDlgrP3Pj5
tFHLEhnDfNngQmpUdABsj4W3EBiMZxunZ/NreUfdlqwAfIM9LC5HN7S0N45cLGKtBlVW260MgvoF
/WYBHPoyOM+Tzif4OVTDmqNoxwazGC0mo1pYWKMoDKSWlR2Zdu6YIy3nw+GaRA/SOCBWMXvBFD4o
9FY2oCHMX5Ki6C8FfPEfIuW+5I9VSelso/mx/CKYbGV9gIo0ll7bjmCp+zSyWieOctdDCeAxh3pt
13Tm36pwMsljMtaoSSpCJaugxldnI2hk7GCE0mjGFZS+P2AE4e6CFVs5Xn5391iLVTHiKJp9f9e6
9C3Ul9yo6kdi46iJe9v3VeDCihEdm39MxiqaI32vE2d5/yVOUCiztDdq36Giofc71KEYUUg1xZQs
yeVn6cOr6QO8TxO6P2XcSpqXTEKm5RceQpIzlHnSiRkHJt7iH7whcVbLpFto7NUy8pC2/F8/ooRy
mRHVfnwXHlSp5Qt9hwm77WKPeZ72szj9YVUwTLebUY1KbYAQ4EjOGmcOWyKgt4+V2O220jQBfKyW
gUzc/CR9Pkys9Y4N5yRpBSTHmVRrVzSancSzy5f6Qaf0Ivr6wfTk6ZG/YVgbqbadBxsb6XDeL6am
UUg2nnRUp9wzDeE2nQOR65U8Zn8nO7LAtlVrn1CfJENLBY1PtR/Ae+PS4BQqnNqwAs9spEm9G5lS
3bKEivB/1dDBC1+xCHKwX/1KGTP+k9Q3K4Z0dBuu+R2wSVz96AVPihFefJ6yTtM2Q/gD9FvuQy7L
0+k93ohytjcT9MSccGWqCVe1psxiUMhR6h1Fk+NN+GI4t1uwwZDWmTWjDSe/yRzNoWjCvBuQ2/cb
SYkyDFkneamHce3SIf62UvDsRROoy8l/Oj4aXjI1B7XeYrYAJ7Wm5U3Dm1ME27hbtJNiUt6OGbtz
UhPp3PFnxUd3dOA2I13nMh7j3hY0BXfhkIpT5+bWRiiRO9I4dd8zMlGLEnOfABFn66W8bIBt5coD
nZotvMsS4bJp3ZE8bot2E2COSbKcejl0QNo5dzI4Sifd3r7W23HJ9WqQawJZjY0vddR3D9suzsDa
qKSV2j/QDQwJ1QvVSMcI/6RrNJynNpIW5JxjvlSI8V9qiNk6PSaDLT2Db5npuzd/K70zNe7KciHR
U+lYjG/8v8apSWEpulv0Nv7oYLCjsuaO5jsvclQ6Rp83rrp2He5hideL/sdGEpa1md/eDggOiN31
I5FYczqbTOOdnzUkhIJ1Kb2yJ/T14Wpq2QuXMvTIEXSFUslxlWuJmjtaUMVA1YabM37ulPxlVSbT
ePz2r+lITzgaf6rt/2yCIdFXw8jO9WNpMRA/cqNuoCTlkUzJw+Gyz40dnhBUN/CkmuW9grEAeVLa
DouoZRk0XGlWm1swyPvE4ihxwLn1A36MMBKz7NpZJ2/wEduLFigOz9AzHL1gLlAlIRaJjUDWspzr
u7CerHvz2iYy07jiTHWADpZx1CNxLC/UeG1uTMDsgiB0t9EFZV947TF0vsITB+m8ylL36h0IadGe
ke5orvTQ7AkUhai2JnyJ4AMc9T7m007z3toX9uRzuV+0PJcI+oBDwioo8jUoB3mSjqsZKqRG20Nq
LxkLiJQOSCN01IDts9d9PihS6cpTk7SR+8yqg79w9JwYN4z8cj6NyD7mC3cvezr2sihiUxMenZ87
xJBCT1XAoLIFzCMjacOQTArjCxNyATUnrD2kIjsKNPwhnnZuDpVzj2bacVSGslfzXoCwynaEIhOu
d4/pUb8/g7gjkWP0VJloD8cpbK+I1g1JWmLXGXN7aEZw5Mig9je1z0TuBh+y/8ZgUEu5M1NpPrFO
2m5i1DH2jIVdDuPRkdFmvmTijDoR6JFDOBubMKKAgTjXrQezkgwJyvj4J6ekOHyUpSzMPH23WHaw
YxCPt4NqhTbGUR3AnXPU5UFhMWRLqj/7/qZf932z9G9qUfm/iIoUIjwoJKdSzBP21g3WXHTM1Xlf
dZuodGHgWU2oXSTm0kUVOjAE1AxNLmlSMXCJFcPj5sX6l0Eau3zd1CR8AJk3IMju1Th7bqnA/GNi
9CwR4A/onP5u+W1fE33rlh7dbw1mp4VmG648+Wx4T1UUssUjUZOBf7CiuEF39jyOQO1ygBLXO2uf
oDjblciYxlmxUED9TbpDw4izchsb6vVMwgNNXGr0z9BFdbNPCtoXzWftLvKkuKRdPKK3v4+fLWnn
2lHlRiUZv/a/+bQS9d/nkd4MTrFyn07t58MflJiuvxQbAr1VnGoSw8nytVK197ltIlJVHR7V1uwj
k1MTNfGl2k0uBtEcBXeikrbwc3X3221gPgh10zwcOQS4aau8JvD/d6H+IY2UAN6HOIg4nrjh5K49
TUAh4GxjRtemsu0DkvyLBlNec21AV37/+4PRCg/WUs9u0jJYfsS6Wmo45JtZ2YgGiwv3tC0HzEPB
/mwdI8zXIs1WEiif2TYDfFfuSQwE66ffFiGzfgDhxSj03LYcEgB8kP+3hXRbqhQ7ByY5FT5CCWx6
YjXhPrdiJor0tByisAV97KPyCLiLlt4Iwk5MLSoqQny4Bv2l0v7C7fBYprVh+XVnPPdOnr1GYbhh
rUbkc7SgIPp7oqNqInYtX9gGhNtAcqA/xasl8a6D+2J36B61c9X5VMSrqylWa9l5GJBGCXvPumzb
OxGEhOQ4BnzBl43WeSd/pJEF/MV9HFvi9CjpD1XfhFYSjunv2CyVqzGFIl4n8K/+zXiuC8gnI02d
cLGwSqEv2QBAvoVm7Hvsg1f418V/u+UqtdfBmBzOlDOpo+gRHFFEyVaIWAtf8kEF/w6LtVNe+f5V
yS9tHrR465z005YpxMyd2wPnUVpsTnBSG7GKH1dbY4lRLdyEKM5Nt8GPW9SVgnQXx7rhvjiSd5CK
W8OnjbkKrDd7s221Y14necFAMTNk1OgeufRjTU8z0tul5s/fDjUBCMnon40TcAi0IQDlEApZY/sl
YXNA/I8NSpz8dLa0nT8H+Qm8VlJ/zA2wMs5mjCy4FXVImD7r8xDpfrV6pjNxAB+hP5E8Q28Q2RND
VRoO69YqMHFAP6Q3MRKivKsNbuNJ4HGWleBOSVlSiPnBQjL6700ouitGMPSCqm6kRux4NCV+6Gzy
pDHw98Mh4TD9EFpLOMHo9WIBkHx0nvSX/g23clKisq78d/U7z/IPeAz8qQT8nIDGS9xTfuUHrYxa
07WS5o1PusLcs+mAP+FG4/3oxKA4vaWj/QbU+fKmOj8TgTGoNWNt9i4bWdh2TnRcLB/PEAQaY4p8
IEfhsrOM5GsMIzjonypLDXSzMc6RZ/nsko2XUoV2XK1Z1Ysfgx6ae3w0idEPQg9Qjp7UwyjlDKaL
rGz/71ZCKAFD9iJdIlLTBmVml7NZp4s3YcmUx/PEdT71IFLltyWJ50tm3PCW+h4Adpbg+wq4vuBP
EeqrxgITJSOM11P5ta8nX0UAIKSjA9ppDXr6O3r/yp/S8GN+vsiaPwbqWzy7wbQ9xkKOFmMCbBUm
+v4Da20kTjeX8W6Xjfe16UAIlrzFAu39KlmJC3ExW+bFAmWDCfujqneDdKEgBbcjdRfm0JCSuTEg
S5mzFxFCw3xXdSkzmHlDF+qx6kCtx8c/LTc6FD3jfax1nxdUg0M7L6aTWCbhyhhAW6hYDfu/SqQ5
smpnobCjTLxtm3RqTy8Sp/eYRH8ZstmYoP+hgsvY6FuT5Z3PHoGmXYHoLa6Qx9bJFFR4jrzVu0GG
mXFxV0uhlC43XDrEqfeuLsGTxHbppMaBVK8kXxPg8dQsdnuJaY97ZUfAduKdnDR3ltV9G/l+bzRi
jAp6L/mH9XeKGKbcZue0IvOgWTZkldsLKHjg7JBBELuTHIB1D8KE1lJGPQSXOs/RkkABK2VrgTUt
0jaWmwpbEoiaYD5eiX9aN6bDTVnQICChIao6CGiBfzd0g7r8B7uFoUgkQrcdiwbxdImfwPqMO/wT
aqGc93Yy5HeQdlHzYi+55fh4FV10xOUmhE74GR3j46vvdz6Q/RbmBZovDSQ7i4bHK94mVdTBZ4Yr
P+jj8STjggqcXiTr8M+PXgicROcxLH86+8DRYqTJA1pmO7YE/T6Rhi09tu01N/Uk8Af9M4xhsACc
LHaN4YyU9wjTbAXPOPU+fA0EqegNKlnOXrYpDbd0UMCgQBboym4h6hjwSufGUAmlt4PbkZqtD/D8
gicCBXYE/OHNY85W1EJHwIhDw3gTL969dhXr9IDEp7hhaFD/SpC3MEMSI5upp6Ad/ethUffBBPfs
HCMPu4xzsl4Vd3bTWucLigE24BKIqjUMZ1r67Vvgq64Itp2jX5JjbLSWpafMCQ5z8lCqOqijv3Z/
p44E43aDcim0ouqonWdsuAsVZzljsIIVoKy1hj6sXMlONIYPr0mjfcBo4FIOLBJrQNmt1fFMx9Rd
SWEo5yt2fOyj/kxutci1Pz64psJWzaNTAYT7yzIe8RHs7VfNvelRigAXKQXlO7uw1JVPPmQH6fHq
x6sDjzJXM5fX+v/LMLDC6NxJ7NgPcgThK4keAkWlqCCGGN/zc9ms/Vt2Yin3X12AvTxVvazv4UhK
vsW8PsYI5MEJaWy3yybAoFt5UTR3u6CZ5JiU//YGaBcBp5+FiWuLAh9gfELMK7ePX6frCv26t2Zr
mx3pfLKRcDZtya2rAIZWs2+0wRjSjsbPL9tBh+dp3+PFoXNLMdP6mMLQ97nLcTTykhohqo0Qemu4
FAI5NMmMyEGSP3Bg1bFNsx3CpgQ8c9LRMXPV1WEV57Gsno0UMWcfzurRCIzjZNZ4VNECQRsw8Y/m
JyrKbv2n9x5jOeWqMCLI/ZSC/1GTPb3WwoV+dVEEbgT8KUSszwQgoTeJRAwYTBqvSEeCxihVjL8i
cc/g22++Ifs+KIt+cmKxJy7hwelBCdRFBH+ZD+f9wNkBU+zrM0f/HRAOuOuv97vs5G+HI7Gd7jDz
dlvvM5gr9AsQf7vErVKjNnKsQ6bH6lF5ADoCX1EvA+/7WhiG9muJ4/YCLmwnuzft6hKbJ7+1Cige
vbwhgrEGjRjlMuBGTCqbx9U3+HemyixqVXzZ0wY7zwbzyITEEDTmOsjEcmEE+gX6pCNily1ir6ci
lK8fwxlhX3nPR4u7xHKV19loyKs1JLmeYWmc+dyIp3vGAq7T2+FvgDeXLPRAq/crb+r5TkPrtOyN
PpPYGJaW8zeXUT09QzDGDFi8Q+c9a+LcJ1qUxHZmxZzmu1H1gKDCpTMnEvYJVhuFmGhcrlviwk4N
5Usdr6+ks8npyL6PNLt4yVWUemvALCTE8LsW+DIepxHiTiunZJVqHLdxecGfSQB4OhDrFNhO57/t
jsoVTeZDHo+5HGOedBmPw1d5Gs+tPs7C71pfxvgZwzSCYtxzt6I54cDwyWUs/2UdBePSdOEx3iGI
ngKoLsj8j6AZWfRygFWuqOW3mNVN+lq5zZERx8MtPSdOuUVXEbYaeRA5W416u5rby0eNo3r38qF/
FeGceCuuTucNKq87jrcpZf4gSnOW83KTnIhsfAo3NcYEHrZprY0XrCC0R5uv9tW6nQ3hRyM1JdmZ
slu/POzMcs/tnCwQnJgeS1SEo4NAiDhN+CVZu89bfE5PQfW+x2zxRDa2TyYT+3C5SqHIeYRbyCUH
DzWV2S0a422w2AcsSYf27hGhtrPflFn/VS3HgdvEKGkIVohRM/IJvdPh5bD66wGTSEn1ycbY/axZ
rR/I683yMSV4y2W+D/Znbssx2MITIjoY1/kFd7BGxzG8aYwYmXX3ROQSweKupih7MQRkg9z4bshN
sOEbEYOllM3BVbG97vw4Mp0OA7e4YHtR3Kwl0BFKlApPirtgiyaVQ2Rb87RJH/XPuiuQSRwEVZ/W
9yvZxx+98gir1bHYrM/VP2aLwT9QHCVLMv++hpCK+1ZNtdqeItByPwtn2INlNGo95X2piaAAzP+I
5BrgRST+VoZY01ao0hubyjb2gbqPV916OoGdWfZIaJp43MRFPnXKQeqITC/4+JgNlhpp9hczJAR4
v5XeDtxFxkWvlBjT8pPCQO9M9HXK1Nhko3t0+gWRnQ0XeyKQwdEXKQBbfLy+i6BZyXiJmTBQHzLt
qdyyDo2MFRGyPvmZztzfgY5zMum5xtEvWTehlGzmEPptNNOgUAHk1Y0pHdibe9Ifj4PxmkTEsulb
islu2wVSCTc+/ppxD17zxZ7PpGCXRCAfxiWSFGBJAh6TewLj/wJxX00l7rZ6tr89LiWrS5rrFTtY
5eq7bDdOHpfyDQPqNdxGJfOJf4F0JlXOWBDyNpd9tIqLw9UaHUSofin5Pae+AvH8FaRz7A9XtKo6
1R3+l6Dce8r90b1UVSo7OhwKwD2HDpN1HGSkhohXnUWzYDpalSsFFYtBSWwLQX5+Fgyqz2504zLH
xZZyjcdIdeyRJQgTP8DsYk5RsI1QO0ZGVNvsKzySZ5FoLfMARIh8liyxezpkNczFc0ti1/bOHRIA
x5YqBMHqxJ4px4Rc7OvYbXpEueSUziTRo8Lrh4GmwFujrE97m/pCUBll1fEMPBpKtx7hSnqBWiEv
o04qlc86n1aE49yeMcOtZBk658kQOAYmW9nhBRCwES7ObGVKh1E/H3arbSvlSK1WOG78GFjMM6KZ
hqQXe+mTk3aayJY5t6PKnZBqB436Kkq/f+LmW5WjZYg+tduEQpfyz1a18SCZiY52MfFkx9ajSsLF
zsdEWhlVfZFmapTirNe78zuTp0nfuVplXl02oMCf9b+rsliQT9XrWQ+IYbamD8p/74c96RuUSYFm
Kl9kZIIN0FRz1PpEZALx5Zt6oaUv6R0SEA07yeHCYlAXeXxlxtSvtqaUH4/11fNAA0cVvMX+jWvl
uBiOQaQHY3l2jZuyvFwH3UxRE8EDhoDql0Tmig7LJo0Jipx93ah8g6kZfFTkQ2DbFJbzbwOae1rj
/MimaCWZ1gtXn+dshl54ImnBeILYJt71FsSiiVO2JCxBlaYMzCWHMdIUphBYW4/tXtiJMfJQuJpS
eJo7QaqUbr5woCims1CvFgAohmQGW57er6QNPjDakrxDxEIUtoKMo8guhFY4WK4b/9E4nb5j8ga9
2iAfs0TJJGITQTj4XPMRG0ahU1V0vcKdUpxe5cVzHry+zZgJ0TmHN90hNhDWApkCaeKtESxf78nV
5IY+XInMoaCA/w1xSg4NOM/IntHFlKMCR/TK/TVkwdAUgyLffbHkd+s2PGqCi1aVyv9wGZ7lPmS+
joW60wqyh1YGOTMMhMmH8cc8MXPQOPpvwIiR1//eR7leTw31RHAPqTj4EWPiHG6YpvIEFyJT1exK
K0dxXDHfeTcfEnd4Eaa1EHCBaq6hbzybnrpFJES7aKRljeGvVcR4qWE9uNN2v7Ynn/vcxLKKags/
u9t8b+i1mdPoqo3NxvY/BJEM3rRTzQPudw2S5wUuIlbI6x/vtB8P8ykSTtR6Al3zI00xmrfWFVAS
GSb/8+1WxjCBXpt1ooanTNLckBq7b0PDJvLZo/oI1VYkCOEEUSdekZCkzRJokQ7lfNw3XJ5YHMvU
qROtVmVyx1Gq+mtYAfpXxLui19Bcg/PfVff7WO+wBrt3X/vNl9FpAOdnfZw+gdbaZ3lglidtuLY1
XdHqPB8CcAtMOdOMrualTh7yf5dFkmTHOq8qP2BPKYoP8dWT/OtKqX/B5vFSxguV6PPknaUIUaUx
0m2J8KSU8eZk+F/uOZI6DohlAft6MxoU5ANnOjhx9L9C+0u8MswrxGHB8ZXnFQ2e6y8zejoHlZat
mW1gZmoAiGd/3SGyfOy+emXY0pyJ54IvDPdZ3GIhyqcWVJohc2fU+ZAnx+sw4yG0xvKOc+qLsAcq
tDVRjs40a8JQUwy/OOc0hco2QsvubExSah3PiPAwIFnhOV42dbgdQEmiraiT2b5jMQO2xPcJ/aly
eyp7Uw+KbR8e0SeUX3wraQ8vxjBTdbVXPw/YLfmgxcf5+nT2274exKj4yB2ZOHT6Gw+qTaku9Irn
uP0thuLpJmgxw6DSrjMb0eKOGZ5snFA+ngp1HgpyirCraSGKF8TJRMg9zhMn1QgDv+/3Kh89ppN4
mH1SiPjpM6B/KnbDdq+kJ9wEB6hJd9xIYDZ+Q2SdvUfqxV5J/ogZUobEc1sCMkuqBAMs9EBFLYy7
EeYe1ZHspV4yOoHMNQU/NCwYE0uDhYOr2p6J6eJV81E0HxwZctb/piW4DJiWyEzuD0aYkPkzXVhy
nWKE42kdVXIjI6rDwVA+MdD1kYSxXTV7Ms9WeiuhOyKQEXf2WzT5ZJU3ipEEIty+djHkDmtweGYU
5X+z4PzCL6RyuPiHxq6EmaiVuOS+Ai7YZIh02nIail0PrMo+OLfHc1VZkQ+fwDeANGSc0Q/q41p7
yXU4jVyTcuO0E6AYQ83Hp4u9225mNE6MLUmf3IQM/y3RPBAje/seFn7GU9ufUKo3uKE6doWxJ4bX
w7FI7git87hqR5yIek+nRdCC7muRVGzWrEYLLehlUfxgWDLdwqI2/dbAlFSrHgtSIhex3SP1oZ9z
lZg6DC6714OP3QBzXtSBCTjY+St4hISCBbNIaVUnSABF4qI3q/4YFSkWAcEajqvmILX3OAq39ueZ
gOEhgl9KJRK9ifvH9+5nhrbF5VyOk2ZVOZtmbCtdDkTiA+yu3W0mjibl9OdI0EtXU/7ZFpg9bHax
ZZacrrn5rz/UY7ggRfM8b4jdzFNC225bjnoviHXeFs74dvuAQVIGYL0yz+lK60IN1eYdUCE+OZKW
qX19LwpjbNfNqaEvo/LzfpsSQJBSW47fKy2AREmnvB6JMjnCw1oX0XGKigBCJcXy4Ulzj2Zz3RDe
dWubMMrvutBXEvRIaRxiqpD89V7AkVHNMLVEMVJ96edwHSfSkXnqoIDsbasJjpSTBdPoApWjwlON
9qhfDDVrL/cLD9MOVrKo16CwuYMbuKmhcvMaSXCiVZ5gxlemVHs7cafIeUzZUnXrH0T5sBPN7LU/
a3mpBKYj7WJWWKQa5KuEupmYNBxok8tpVP35gmC5QQNM1INBV8r3jYuSXZ/bxtDKjYPRQzihiqMf
7q5jZDMJ/MY3eRr5WvtM4z6BxleHTdoSx+r2EQnLP4l3TrV/XpImA9h0T9+JrXJRdL4Yq+788v9l
a+KS8Jv4pc3K1LYyr5bTJAkkMnWI/nucWSFtNInwu/GGGrrUPc6bIdzO8xw150Du6lDcIj+e22Ml
sFjaZf2DP7SfDZozV1xsgkGo/nkXQJQ3WqvYOqpyRBl6PywQbxQyeNzvGOpQzO43/11tPRdgxOAr
imFpf9YXeVY/U8atZrApFGrviVYF4/kdM98SZu1akDw+RoByMKKQ2A7ixp/UxOMHThRXXeY2JDkH
eZriVfj7f7YPgRsK8MY+6t1zevgKyGAEuk7jw92tPVYCiSZ36uq5pW9QDLtmV5AWPNT3ry/Rsh5E
35rYrN48oYlUQFEbSupr9Ny2RzUs0od5OTdxM/7Wxn6iHGow/EQVvzaXiNiXCqbhoItrd+v730a/
seRnC77E3AFlLr/HDAxd4rAF/6DZs32x2W46WhBjMA3T32EJ7FnDD6eu39liwBB3tZC1qLfZa1Gn
lVLj15GAqNc0UJWrRGntRGB+iBi+e0UNo1tV7knqYN41sZbhZ+bqNt/qicIRYpST9gH9C20sfmOm
d8IETxnBgXLkTUJuhOFJayWkRnOH1lA1l6EQLt6SkFNu7zuavQrRYa5jjzBJRpWelqY2KsY7pMpG
I22LOjgP2D/AcFK+uBls6s4xGajVRa03ZBW7A4o/ZQCFTmuE6VyR0d1lpugefPLJRDooSV+nwO/r
8Id4P9v3oMLWz1bbW8V0ltJxwE49DT5Kg/b/fgsDjmKTu3L0jHFgqqXOSntfSS1gBULNRri2CQN9
4jDZpG1AMiX/HzxbvPj2o7Cw2A0gWSavQUzr41v26HuddNB3XWijMrh2ECwMFTK97oxn2+on2neQ
Z4YlPWT2CsIpBgCI+kHlugXqTuTSQhmVDkSB1/hex/zlGXo1JtaG0xXFad6X8TJUC/EVZ1M0+ZzI
O47HN7ADJ1yxx+zDlVVKRrQxvpAvQa/xjjQc0Ozp4Goeygyj+srNQEe97/qSrVAo6wHgZ/L6OfNH
vNKU5aSYdOI/a5zuwAemHkUqIi3xWJn3TGLILXSaCdkyr0kid9LJ+k/xYbQRfkg3zrXZdfx7e3dE
hc80T+hXXgHk8vlVslZR04uxcLWVKm7YXmcnHF8UgfdWqN7nPEfDmrp9WvnnqHLf1YwCHSpZLgAB
7PZBoceYvuxEZ5FANm+7NbqTMSj/sJFHbnCBCZLnijGcmz265WvcSYEgbY13YoY8avU+WpT2/oV8
cOf9oWKKIDuVKH4yCth1/aGtl9ZhVp/6etDrz876rsw3DVWL/wW0Cy7M/AckbMeryRIQfAlmkUzv
GYrCvzDVMOf4cOy048NeJ2xnh1ZnOj3bSZv6RndJtbZ57Sr635FpHIrpUsDUKwg4Mk6pwjY/nLNC
tl9WXjDHe/Fih6OQmMYRvgJxJFKUpNP3IJ9GkUaHDbfQSq7Cc64g8yOJkh12uiidOHhcTnZ7EJ84
8+zbA6RI4yeobTmg1sZK/vuTLXhS2P0rmqn6l7pYTlGyqEhudzlRQY/LkS19YmqaCFRftGUy6Psj
5rtURs00xfcYnVnK+fqf5XzeZO3vjp95JlLMB5U2lsYZhdFteIm5Vk139Sht7WKZv9Y5678KL2AG
n4bTKG4ZMB/6hLV3HOk9m0C9DfwflPU3oRc0DGBrIeNfrFnrYkBoae2vZzL5rrVsYGo19N9nq51Z
PNvpeXxJZpJXvVh515qYByDadIcL1/LWXTqidqhKwSEMLwEhyEP+GOnzmV0NO27PD4gkdyCoL1XL
B9X0X0ISa4JoEvi0uVJW+EBrZFUW+zyvbBIs4LuSZI9V7XuaDji1x4OGB4Oak8PoH0suqIpnpscA
eOqcQB4V9BGFhzc2mkjYRLiziDNy5XyFK4tcccOQATOg6Zssq4jSbMOcl3a0JjvRD8O9heZ9ZOB2
WY1TjqLLB7Fdtbjnc2rhbL9qmF55zxQeN/uw1yeE/YDZFxnI8ajz64kY2OCKSuRyNTQy+CELnYEf
XmxOQieiDQAP/IhZdC/osM/vn7GL7UjcCj9tY9ZTwlf3A5x1oxJODpuAN64n9BpOem3+LzjScbBV
dWu24ZIMQtL3T/2kvwv398HiOorbstX9mbaCEPFZaJ5zAN9MF3+ZNvkvg2GzQDS+GwJ7e56eqLIm
ShDH7jqQ27hWwBO1LlbcVsolug1wkI9nAZqdp89/JZqRMGseE0S/Wjs4daHak/At0mMkTPDq8J8y
5gMfUNykZTndR2aA7rOHb0bKdRwXtcX50XJpWPxfjoaXC7MTOSwVQCp5T+2cLZ9pmq1WvqT97vWI
D8x8hn4QdOEbSKzYK/YwX3CKMyJZkWCf4T3ZJ+BglEzBkgTnmyo5a2OGWSrvhIFqb43zp8wtJP6B
tnhdy5nuGc6k4oabChS6bMg1ptWvaub4iawFr0JTkRRpVPmK79Cv1ZwQ+PcupANK8xCV5gmZSkHk
D09oyo+NhJtCk5UiRyKlQucp264DLsYxNP3U5B5bn1wPdfEvvFiE822ac7PDopr2DeinNhnHxr3V
QvX79O47lstn/Ky071bTXrLFOIHVtCN1QvpZZ00ErIiDhxQGlaOzffXFiv4KSsW7w1xBuz5wdwog
QyjF9ubrx8t7czeihZ2XelNjQg+LAvNnCo/EnmwQqSwPgcnyTuORuu4A3kttvimCp5H2/F8w2SIg
QSWiH6Q8/jhUz64ES4cMEOGzrhg2rU29wgkjwW8Dvwk21KlNJLDoluojz9GO2IQgriF/bOqiSBlC
IN4mDBsMnW109y46CJ0YcDA+1nJepcIa52HS65Ahj+uLAsSXfJLJRhPgKJzMbrDuL0mBajdkJg+t
gyhjRO1Yd/GWxUac51MsP8y2PT4gJ1aTFQnVYDcm2ii+r7fCZkNtbNaQJ5XYvwB7+gD0AqEb+MtX
On+23w05tso3LtvikfehknVB1/sLkG4oB4VRLD0Ua1fytoO3CNJ4L9I47rIj7Sd/FUH0asMPydCN
DLyh6AxF5sRYHZ8ejZXD0QwDsm+uAotWguSiCla1lGykSX1ilX+u9XovgxMEHFaNFB0TAnEhGLnS
z6oAPx9DPSQNIcG25XAYJeTASmYh/A7rRZOnrEIA74Wrx2xwQiCi/EMDKQs2Hv/ixFKzFuI8gh+Y
5Rcr7+rxoBj8HOH/Ll8HGAacNqbmb5TjDveLmmNq+6OV80ldkI/cJTvrm7EmpcI+Qm0OVzb2O4EW
M3yM19Q3WySLXWUlLOv/3a0cke4UlJihAmlnz/SUy9C8EZj7GObxgw29uHSGUKZuIeAXUqsAHcIW
LkUGhtlWLV2WNoKFv1uaOHr+LacKw0ejnYImlx6rn96whmn4Hg8/QLA2l8cKXPCG4G5yf5tsqKhs
L7+1XqY1X8vfB7G0CBRU9oQm2GtmH3+mj0Cu0Kjdf4f2jdAZPynMSqg4wHoQIZNmNi1JKnIeAG9p
+mujJAv9hGnhyTii0+CCwwaPS8YRxpL0LADrUx8focLp5XqE4qETGrbb/gI5Wb8zlca2JY9wMUIZ
0/D3MPCQw3egx3ycl0rCjL7kuKe3ADHW38W/nBssL1TnHHA8jBiK9XFhTC6Oy018aXNxW46S13I2
OpY6M0HErswGScswOwWMJh6oLY0ZXBOhCTFkA0nNk6oiaxg7KXcNKRv9hVTCD4xdcj6L+uOrD+aJ
FFMdiMiN7vuEL6AgPZaJVZ9YPh0i+GGrNyve/1v4MKiUv2Fmzhc2GBZMGwDwr2oP+jIJDGQN9Tb2
wlgwRQgESc5P/+etSS9CckJIMJ0lHuv0uW8NjWf4c9Hw43xMejIWGTxho2A8TfiwzQIGNKoAbAVj
HdQcD5PN2sJyqUFY2yTAH7TAbK2/c7++ahevjWbANPargHQpiXMrTMmBOt+dd5dJQSxHDfSTJ6WB
UDpZnTM8y5zOKcCAE/VNlPsovjFe+wQ8CteoGMNzXlbCz4p+FqbEQp9WfvyA58gVEMoyuznsIYbz
6eWoVoTa4g1BHYWPHpt3948ps04L+oI3KuamVXMyfExqWHBQ8G6t+MfrwSsprzQb7nyVMiSLXZ7a
YhGlLFPj9IIrwfQDP1+8pGPVkLyamfE+ohZtJNay7eIihNgL8K3LpJ9yF2J1kxwXXQK2vp1dV/68
Nk59J0zzsljyNtKcJmWYj4Fu+ZTaH3Y8ocDQiaftPge/LEitqdG4Ga0+M8p6kGLkXXo4nNVdG+C2
5NQzFxMDbieZaeT96ia70g5UI4jogiFG5r4ydMNy1UYp/+McLmluA8LjOikNgoCzxWI7lfEN22T0
RshsH+Mcv12+eRFydwYoENhXJO6All2TUBD4FqDRiU8D1ijR0m0keSW1VE6KBSUOSe0OAph8o5xk
2lma097WzSIvrlPoB4ev5QDjPYQyJoMZjvE4uspfZIcCYxB71wgFM4akb/8UIO2p/vk/R2o5wzzz
nC6o17Ajj3eQ/AglSD3V/KPT+shZ4ppPac2y56rRjSA1hG2NIC+pSH6JFMG2AGh2x3BOFKGX9nZh
jMjdO8Ac6EW/O6UK/COudQFF3lCRkJZIc8055cgJTPdeJoBQ3WNRQK/y4hJlUaQD+HMQ5Dmwsias
8o5n6UGozBGg6vsp6Eeq3PjrrCVwynsZ0Q54zQTHU2aHrVeE0oYD3/kQuby6ugbJj2vdIVXTKjZP
fvol+vdR/445KFS1/yiCTdjUzNsc5ZuEoOegJcfCivT861XWy/OYLxUNgt1hJJXLk62pg4o+VFMT
5CMq1X1XEHqgvNnZodwiXloyXGvTgHLvMJ4VCvEvm5IcGu6R5PnfEUIeCqqNmjwIt2UGgunc3GBO
BApr3o8i+VhXS/VmIww6/i7D8RRnyX/7p/vQCWL7aD+3xhUMCsyh++BV0np9OTTQubxIXUBtyT1C
89srTOzzP8EY88964/ghJ5Uslw5x+eMe+SIoQ8CUPUhsqn+BOXd+Vpo/mvUnIB0Ne7biqbJRXrjx
7qiWDrFbFInFL8knIoVVybIBqGxsjD6WxF8vQ1/MM/MIfeiyTy4jrmYefxXjU09qqW+KQ3QZcnqZ
E8Ry+HRq7kdNTbAhv4XdZarFG+xFGJp5mIezKgOivrOoWElOba5ps3Dg8RrEf+RQv3YsgOSfEZGV
KxdeRzboPamL1bXWye+PMLTY81v/+VU30MK0NmDajE+dhHTsclB5Wah8gSTIqEdB2k9CZOCpX2OZ
Z6tEUII7pnKOZQMw3n181eIKthkUj0nyBjT/rJOQmXGhlFGxQ4I9PGsm6FAmBYz4vitqUPrBV59J
RihDLeAeNPwQqdqDXiXFjKgfqb8DprD7eri6e7jR/kUR5yZygzRUpY9i5alq2BeN4yVz0nS7Vxzs
SGyYts9Mt9g30jJvy5bafjstQic0kQ3VCBIcPlr7xEMwjOM95LRCf72SrDn359Fc8ISZ5HgqNKC5
gHA5Po4QYqpGXPuhTOZL5ANL5dgUzW/5Uc7e0EZIn6q3DGh//RQSQSNEEYLX4vYXqkKdha6kVRuG
af5jkmnJoXbjcohpuOpw6RYiPGMaBo86chY7JBLNoZz39XjMx/WUNCRkmBB8q2h7V3Rn74jZA9FE
DHwS4tpnZuRQDnetffrpeMyz8KtBbwzbR7KAhGdoaMh9kK7UAWPZGiy11Ar4m1ZKYiVWMrP/Eg6f
9+rgjMFU1xxvSq4EDpZiuwNbz9TdTExhMFWwdOTJQhUxge8/ZIo9lbhcGd+WmU5Q03Qxnk26/YgD
yZ/96Hwi01mhyOqWBqpud7B22m4tmklZDAmU3ReXxbKGTt+mW9a/YSf28oppiJG29Bhe5o2Z55Eg
1Fj2bZBvDJCY4FzMrWXa2QH4ZgOHmjine+BPROg9mo6ngyAPtn8z4SeWhOaAt98EpjX6A3DnR/sB
YDF6dkvyhQjjOATgVLpCDW82T1LywsMasVogRR8iQ8ecghbL5SaZ/tSmZXJflrM1WOqdG+oUW+N5
5DyZHIir4miyuJCQjULaQUPgpU3XpkBe0bUSJE8jNM5AbUrFQOA8Yzn49aOEbWepJmmefF48aaER
Xqeid5XWpsAKJb1qo4/S4vUOaMUPnMjT70og8HRTJC2MPS5Hxrv7+2aQGd6/dWq+VD2laXyHuOGa
gHqMGHuWuRUeUDWSnIrAFVa7I97pA+iasoIDHEY2uxsOKklCQVIhwrICjdEvpKAysB+xD3wKRh4k
0SQB+tNue/qYuZJUK+TkjbLY2VqIMOasZeQCK4YNmx43603MaOnt5xZK3k0cbSLI7gKIgLIDpsfB
3OdCr8d3x54wpKOqslVDIuNb89+/0o75NRPfUJxm2SqgqwH2qJEt/pz6FPqQOSh2KmZjkA8fBS0v
S633mW1dYiqe7VW1o3ancr5UY522cXvntHnBW/qyqKo6rCN3UE0iR3Bk4Lodf2ZjR8OVNDUYIkYI
pI3GzUPZzJTgY2kQcrB9DCeP6BZiQ6sIOjMxwjs2I1qnNcF28JRQM1ufZzxNxAEzw6pHkMMp0dz9
ag5hsoMiHxC3k/l92KrqXtwVpXswdh+JIG9fOHDDCL+WN2b+mrxLLvBOI0Nc3hPWbpAOnaE7f0tG
MhUwrtZck4k9y0qz8oCYDexuTM6bfPzzRnc3RApBaCnMIOjp3ID3QUhb1j0aP0xBLh0U0lgie/bK
Fj7mkF46qVjGz6lprtYHOMlqeZ4Ogd3MIXHbS7munWmZEiTOW2l4MySCqyMm6jlHdcPDaKk86sNZ
YVtkBkdJBCWvp4iNuwnJ/axVIYIvHIakB/GO8dwBwmbiiV0eaBzv4JND2AuMAvMnlIUHvnS/W7bU
Nahx1PGIZJ/mTXH0ZaLzdX8BZBQJMymZsffItw/LZEo4rxl7y2c4hhljkGI7qjWWlh9mpOkuXgsY
Oao7VgjjO3Kx7fvZiQRFlyeCMQ392eJuALAQhG3wtCQP4sRMrp7qYhjshv75wWhLQKVXjHYaf0K1
EF0mOgD77jCvEEGAiubHJHuza7SX0uJT8dUAJa5pVQQuEl9E9z8u7MEu51ylF4hQ5R1TPk5nNrqe
uVRpJ38OKrt4+RKTRHK/4CZP2UoIxtpT7lAllGP1h/kus4ZQe+t/5upt/oyF2XLTwq4heSmR1B2S
j1Jm9DZrznYpAdvIPk7KN/BAjg863i969efSXCe1P2gqnwqQgqPd2gpqrIlG+rxmg2SNRHBQm87N
valb6KZXhw2V72mBV2v6dlbEP3X5dd9gXgSuv4vVlyrZbrlDen0OuzdTDkBMU8M/kV8Je61d7YVL
RlYgOFdmFh2y4VTrimNyW7ft9p2mj6uEcC/6bzQ6r01GX6HzwcYUXa+UzjTZDz3RJJJnWULpbYuB
4nae24R2A7YxruLiIMkPijRV4NkH4b2aMHF7229uWLybkbo/GyN0z7shEeBr15rHJMYaVpeP920C
yaiv3yXhtSqnr3L+fovrwFf/puYaBwTNFW9OrRm8EPNRNZKrJ4uwawxQx4nSooes8c0MeYCygg4z
7Pdb5imNtGL5HDikj8F/pRApVfGdixy+cz2rwDX0aJO4GKZWd/9knNEkNCH03Nse3rFc/KU8W/oi
DgmltuCOzmW1WIvZSlu+/3lSZFNTKkyrTjlbJJI47FDcaGxrWHQp7w6dJ+Wt2H1JJj3T2GT72tpA
20uk7/8IKVrglKWavy0Ga6AYVIE60SR+De9GVMVl0ZI7+Z6W+BJdNz2fsAV5FeSZanFLEdX64nqI
OicoJoPromhkx/R58SXFk3R/olWfdqGX9tbG2aEn9PwXorjJlkV82zQQg4QuQxXjfz3z00l5IkdQ
gfzL8b0qac7PQVLF/Rv5FTBM8KBWjytGt1DM4D8vpcIDP/oHHhSlMZ7GOuxHyZkVCVdHelPsX/IB
sAnsEgwAKl3wWMbg7IOBO+iYwVS/o/78A97veKjCoS1SR2O7iQLcHTsOtHJmzY2YIR7VThInBCfU
1yxTXWfHONq9XGkOZrnHvQnOt5ZQOOIEzIl3eLvfR/mKYgzGXXRE+IUbhD+H49DMUW0A0d8If7gF
PRYCSWxVDvsJMoVk6iR/yI53aEyHKYAdadjd3D5GbXDvm5fo8/YsOCB693b8VfQCMPIqCIan58w1
HgZJgkx2AbgKj9zMHDcfIeHpbrQBJMDH53K5XKx62QtIHvhvfStPvXIdie5xuidlYKRkTsszM3GW
p/FedvaazXXskwLLmfyxzobJDPydH1zux3qAsac44mLQlFMAzpgI1PhuvNrHrqfydAUOrL9SkV8Y
CXQcxAJ1EMPE6zLKqDjnjMCLPnzVY52jSkA7Bnnkh4Q073Vs4kqEmdcm8q3G++DYOA0fjTLtZsop
HEzc90Bc2WJ20Isgc5mHFjF7ZjGLo1IbGKckryrC7cnsxriCXhav9pY8DG6gRtzyI/zRy+htiOKU
ibhxSUsFjnOFTb8rNpODeuseTNUPhLX+vxs0B28xGtaZ+1dGc/z+wK0ZpeTG3Ch7Lhm/VwDF0MHU
gZUTGvdNfN4hEuG9dIIcEtuL8Gu/Ib4paMtUsR78hBIRgP1FFGUxpKMB2rgfeB/V1GBcm1v7xTmp
RNqQWnK9QZvhggjjLooe2+gLdTT1NP9CY9pU9KWpBkb8E5ku31M6zhVvFbk7d0I768E+bexMVih8
qf9766nmIDr+4RHX7FXOIFefnuECVJO2qJKQ0y+KbOHFZ0kKh90odUccLucA1lV5KI1Brh2pWSLN
cpVY2IfGXQA6eMluzCM9wECh0kYrEam2DUcSKw/g52kR0RYoJdPYjFiYmF6RxnCyVGuOPVq7dl1G
AkzV9naAnTesNu+u7TH1yNFEQ4uXpb3DvEAHc7ytS7RECkVH5jdEZiPQUxE+LJOyGG5v7hYt0plP
qSdP52eOSXxN1Sk69BH1by+x5gw+GhuKfBDuIVyvXL/Zbz0HrpcS4VcPO3iOwR8m+varMP/jrhYu
BnmM5GJaUDz86Vjsxl8jQC+k2oOsaNO5PWKV7y5PdJRAKmpHb6WLWDPPkuj0GKEFsliauba+bEFl
GtIU7cu4RGOEsdCTEaR842GHhVwnCFKp5zTc6njsUU+fGIzlTxyhDxkvGvq/FRYJdRkP2AQAku8d
KtKWo5m7fI4jiozj9ul/tXHWU9Q3VWsVuahTfFPRXEjaRb9pxWLIUJHc3eA6dVE7zfS2lp5+CrGv
S3vPX5sCCUvp9zqPLrYi72OBzRYg6kmspdnIwpQRs6NKXSgWQVBCOKtG0yu+66fNowBmeqhLH5c2
xCVyebriJGggAQPko6hiKMWeymfliVDcv9k7n0M83TWNkxnY4sJ9Xj24fakuW5Lfg1ZvjymOiRmh
7WSQD1C7jybznXwEMEjqrclLxWiu/UKMZk2mWSbnvgB+JVQGpi0P6fvWBNZhc+deWcbVQkE1WRgW
8O5A3HsSpxXdw8iicoUKVH1SNzUNSTojzyM+b4xPNTPWMvIK8GoVoSwjnS4rwYi7HyUq1dzlhxxF
+vGrYODvKS5Ie3Y3qJ6p2s3YcT3ZqA7QFq9AT6+1k/ETY010ksyll1Kiqhh6F1eX6WBKJKnQCneu
7oIFR2WDhCuonLEqF3tlH6YQJp5WCq2iOgHd54SoM1dsFYVR1mqPqF3lsW6pKZFDxSBykgWNT9id
0eB36vZ6OmrOGBMdDeQysaYjgxda/VUTmVz3TYZ/q8vXY4zhEdoSjsHA13GJor8dI46s0bVKOJti
cBVdXP1UcSgAwTVPJj6+3w4j81YG0MGDhG2NqgTrlbnDCCtQjVJVhCljH/Gky9ItBk63YTJ65FdQ
L3i8DnX71ORBcUb9RAfIxUt6ajHD//qAOFIMrQ3gbCCNVmwW+4bhxlXjVAEkzga3rmrWiXxNVlT/
bmB0vbDH3pbWGtDjFXRBlSYalVJl8SR4pTh18a4Zh1TBeT7178L9lw66CyMYele1ne+y3tLEEqgE
zJa6AH/FKnUe3jHQoEg1GP9LsCXWcGP6fXBA+yq+J9D4mUDUXm4TVXEArsxadIYnTI+sfwXjhXHD
U4uzNv02Cf3FjTv0eupW42W4dboypR1qzGb/AN37Aj0EMTsM7o3MUg1YDSnp50M2QMEi78ePauNT
uaVbRx0w/RWUnaC6GSH3VnsYZB8exemkwkKw5nn1ug01LYqGkyTkiDziGr+5vAUqFZ0ou/gc8yZo
LRR7hWqO8qTO9+wUgVjUfFpwQQI9RVxqHh/QzpxLxEvN35aDMDCqxwCy0QpbXUhmwWzg8z06ZTSd
9jPPHjSRWHSlOL0sG/BIJuFbLWJW4PXRpiRva10DsVXfmIRSaUSPi03scrqaj9gpvh2SrXxhQ1+P
hRgehXuWwlWzzrR3LpOl88aAJe0S3ZPQ0AvqTqyggUHmQw4F3QznEKEiy0r35OisCNXttWx37IUP
DU2m42yL6FOMVG2lB2KcQYoj7kexrpPs8lpbrId3EhSN8YxLxRoMfshaG61Y9lzL1aZxZTwVwwli
deA+EYPgggh/kMTCsdXI/XmkKNHpynqyErKxYmYmVVxeGOwWjvuia4pkk0815YExRLEdMIrdJvBH
zWv+fTrxkBUwwc99P4UaR9TGlQ1cuirYhO3ogEaKb/5t+jAPOE97XCNFbryZYk3UvqiANgSV+3RA
igO1qqPVBEYSv+7nxfl19FB28fbr9TvUyB8WS3uT5RUydJXtMJ1QxreL/12wnouqqYWt8TVV3PiJ
cxP5ckHh5oX93zGppI/2IiSQ1UbcVtpNs0r1i/8bWB0ZJppjSvYgGEUGMhtvPoScXHfTc9zREPWv
3qfEdU7h3blNGVsO4R7NVVH9XTiYVv+V+FwL/6GZxmjV1Pg0Mo9mhXUXVUvmwMvYzW7msyX0V1wJ
gL2MMwLW5zxDyw+As0I746F42UzZ1+cfvMKQ/HLQASX6kQrjfP9b+BoU+YTFVl7Vqz7KkHbINFBp
ZxIDXj3CTNZc9DRCOkaeGq5OZ36h9HO1Bg69S4q9+juCstHZzbOkfhuYgx61ukGg/BuC5Xyln2RP
jpRz2GAbTZgzQn5dRSUYYRHtX1Lz4iZLVK26uaHWFRPGj/CdrJCGeaOmrEWPcLlNSBptHCwOmRYK
R2UNoUa1AQFyUMuPUMpU2lH8wKRxd6Ggnv4HjRhLJNZl11KMAc0xb32OaypP2mn+vK8l7I8oqT98
rcLrtpVvMuLzw2W4E+IbyTqX8TsCXnFT6fjTybyW6QfFA1DSQ1XUfhKGZkOZ7xsctMRP2W3UGAB5
i1Ou75om8oGTd+IUxKYFS/EeTNz1Y9s+OUCT+eHCKh8Sd/B4dg8C7UAgA7XuRFPEljGaTGjZD2qt
Hf6P70LH/SY1igfMSyYwQwqsv6SiIlOw/rlIcXcdhRwmz+P5govg9za5/uRixPPvxUFcRTKWfUWS
+vFQXtS+pUFeIcgAe6FFGoHczvKbi7J/5PPC2qk8Q8gnyvY/hVYZ6Y5WRq3zaQ59DDkrvsW8/gSU
w0NBcmhD+aKqOdDlfu2gqU9KwaVRgtyjtaxDaTTlmkFFQaQM49T65/S0cUHHDAEdo25BdebhAdJt
9f/ot454XwMw8iiLAqV+NsRGWMcOTe66zmwpx4tRWL9eAlW8R/rE31AIPoh+GVx/mIsxpbz6YO+Y
RjLiptNAhxa+wrJej8izY0Z4NKvnCmSyAktTAgNg88cMPbuEu0m0cG1olz9KEMRpSljzt6FlPRT8
WopupnFAH5O9h3tggX16QT0K6AEolrjC7nSaq3LUjqReqzTV6c+Dvt3h/Bgwbcvid+Y3Lqoel1rf
MgE7t08rtXT8AZ4sou1CMVpzDKe/JzUVg7GjKDYc73Nez74bRoZ6OS66BAko22hIUQ07GvPZX4JZ
7enbNFQTx4ok/ajoywTgXAFCl3b0Q2uFBhoFkI260emXH0xuDyDTbBIe6KF4vMZffhzYqDdFyXak
KcOLMe7ac+qtQfHIDUWWA6X+NTCDYHTwGUWmAnzlY2kqtSpfGEsuqtdVWk2eTf7k+14IWPsehVWe
vZEULR4UVpJWva4oet74YbcpEuzpm+VVUyaEWW1qZ3vP65SAV3A+HoSO/04eX+D3pKAVsnK6K2BO
FBVmLpw7uFGvWDPI15EJx2XaDwVjez2yBj7Ba70YZXv36LApDaW/u10E7Z1K/hs1QsBl+o7wipZB
WuKkwdl4yXTDPJ28qcygYYIqBJOReVneQsDCfLh1ihTbMIZvEHURHEVulzqBF5rHn75U1UVme77e
OJf998CPLpnFDyJdSe1bcGsHTTwTSmy0hOYJQ1qd3+r4cEYZNhmSjOWQTsSgJ7ZWA2VirZOuea7b
uBliEbkIE5W6GuzUe3ivYjPwP8RTlGVGsFDGiQwEB9fu+rsk+nVt1k6GZhxQDSKoAW6HBgdOAji2
/JkU0keowBhyyp1NkZ+AX1fDD6xBlcUsZGjC1ds4zDhcnsYYOl80AZ0lSXD6MNLjAFdwFt5cdaeo
8lES4Z7+dHGKpUsQpK0BSWE+aotZbgC6XBJXAuW1oEvFHHN4T/2zxdvIG/9F+HuphhI5VqvU2m73
FFR8BZAGBH3W/HDtfq5wu0SS6SO3uSjvfHkslrhza0OYrZGOxfSwtxd5dwzKHfCoEtgHvVO1+IyG
W8VqEshSPFoQ3z1/qJ+dYM1LJmjuj1pMnBRa11xiZEd/6CekCeuqGdfK1j13yzNYdfEQWzkPtbfC
nDRoVQDPXDM4psnT+0VHiB9I1gAPoTYeXjPYt31ki2Iym/Mkhv67raaEzw0q5iJPVbtFDSY4nyIR
4kni+WTvf018jcsrF3yd1E91INxjCtLkqu5L+axFoGC8LbFRaimnUzPdHsVzf47jhumrRJKYI07+
SdAQo1/05QVf0ZsWNd0QI3oTwIwh8bpLjk5OhKxaBylq3XJa11umYF0m2asNemU0+06LB1UbNvWc
q3xOD/xdOtu+vY/OwWxEvfj56FQSHdG40Jnjtz8gfVRGyfQdh4Ge+9mX/+EhtezR+loT1Vpj8yD0
3y5+44RM7KhfdEvDeAWNVHuWa7p/3J4JOxYJKzeitjwpfumJO/n4eGAG7n3FTE2I5ZzrCSr7m76V
Oox87pMUul6qYp3Co4X3C+bKmKLdugz0jb8PS5Ovut/ySRYJXNGR4HM6bVXrsNM1g7f4OTABIC/o
ktzsA0JCZnxsPvZR4u/EUxAO6uxOFCEKoD4eMXlYo1cHUcSunV94EHViNP+o+Z+bFulRvFPKv+WJ
vi06oqRp5EHE8C3H7SIMRPQcaEbpZjI1FFxrwPy4SqTISFtzvekhy25On3qWRLpqeRDY1reYVIUa
64911+pz7fNRUAB028jZa8MFCtOoME5efPpI9HjK9YF2sBJ9v3UpzUAIq4rUBXTyNMNtiOJGBYXV
uNRiXe6s0Po/20uSr5+UrQOci3vV3D106BtzjE7OYWzrPJIeVMoAJ1VaB4ZHdzWpjinwJl+Ys2zK
NdRGVHsSAV8SaExIVIdwZLkNQBIxPs/Xnq1/ZqN01fHtUKqCX3kxKxrmNaUuQHDkUI+NAsSptJbY
almYkVie6ugWaByKnMSZMdwDigtE6Hx+hf0/5DQ/XarqwAyKwz1fhxJ1CcjOIcQwI1Tu+TyudOgy
sNy/8SuYNWlZ5RBaGW+tddmbW0SEawNpnyKHOFMEDXHwD0haiWs+R3XGy7+NfOsmrv7uVXgiBwXR
Ojde79HwCvQYZybNkJ2CwQzz4PRnLLShYg0qFbdWKSS/3TjJWsBXKT1MG0X3TYBJ+SLLpJdEjjLZ
jg7+8x7/xGbIHQnJvjUblyGe8hHzemsnmpgSx3jC+pd3IwsyfMKkZee1DTFBNICpcdLPoXGLju7h
3Nye8YJZ7BSSzZJZF+9uQ/YxHXS6smg5o3jcOWM2YjMRCs2du1TsiViTfFKMis0uH/JgTvzsZLA2
eQnfi4YugvGQAC5WeDn46nlnGkZCJmmYMA9erp+70I+3FCGr9u5majW1C1LwXQpfq2WtwQHCqi88
vbmDOyXT6sTHWufGIHJ63oftXxzHUjHT1wODV6Ab9J8Nc8DRB2bWmjz+L6w2/us5B/mE5nX/LYa5
6CXQKLmNEKouiYk2sl/JuTO5ED77RsiTsGwcBXJdpgLuznFaDPVxHdzJw9vLczm64/jN1aGX2wD8
5snv+jfHozd3mdEebe6RlKeQrOR9P9bot0mM5I0gw4dfFA35HUBmTYUiupA1RK7AXsxuSk5NSmOV
ILG2AfT4VDpgRAkem5NGWWEQeiB0RTFDrYo5Z32muHHHyb+nkAiTbf61MIaJ0/BYLdMAWciceSkG
0Vu9KFKhzdYMBh1ilhSiQzUmBIYOMxB4/QJ70sQp8iM/GXP4JaLIJrBzl68W77UB3aiDOYxyFUUE
IrY2uERjVWRFndQc7L1ndWahmq7lzTJ0E8PLoIuD4MdJ85+ekY7BEbevopxn74TrCf3VSYfeuKnb
qyFtDjAeMqt56yAb7ikfUKTmy8pK/bOwOAfy1cI7JMOuRtwVsn6kU9TCzSSzkNRt/imT+V/WLYaK
C05REehC9Tt8b2D82rvBOaQ+D1j+tvrtu4sbXEQB5RmGS9zh7ZLeKWc/JbhJFylUYLO+MswgBTul
O0cFzhus/PD/ebfxLXKHrsUOI75kGkUopVh62eOZKuVsKoM5mCLHwtcZ1m4koJwFdQ56+UykgO7G
RiNMc9gzuq2CkD+Y7/MEnDd1/y9l0UTzKSUbJpUl9sT9c8IHA4sMAaYJsnRzM0lZnjQOPoGRsI4d
8cP9Z5HjoggLi5k+CpWjUCt7ELzBCdDdT205XXau2WnZb/K6MQwCBIKVLGWlIjerWfaioqD9nWjM
hbTacGpMtF4guW1FssguIYTz1B9H/9YyhuIWNI+ltEeyDQ0f7TmR4cNo6uuTskRD0/E+x7WaztHW
OGMH07VS7DZLFCUVpSAzL6r2OjTc08uvx+BZfj5pGV210ctmitPiSd3LYsP8M9zt/9Qz/l/MSkta
LGt80+TAxAxw9IT5rl5W+uHoTPnoroFfUovbJvxyok1PKJ/WohccLjoZ6dIpLpMfVJV1aqd+bGr+
MFH1I8ogB8EMciP09kEdgAWkO2E4q15zmBS/wuUkSiuHKfqb0jBintIUBH7C9sdr6K1165ztZsf+
6F+TNcZFuyAeCcWvZrZU65X/ngOO7Tr1pmWOnYicSy4h0v/P1a4BP05+a4Doh1/QnMLjaUmDlQfa
JcXx+YB+i7sDo9yPZwJut+BvaygRkPWUX1Cmh/s0xj5jogy0lQurRKaOdkSSRb89PNWI3uBoH1ok
MxeB3CQjFyH760MRmXbSfmyDRwXQNRgIs1l0kqxsNhvrqScOf1jEUrqhISuTU+AtN/UyF2z76ef2
FTGLA37d0axt2YkGQgBL+gN04Uhx+2zl+/hSW4azD65IC8XZdDQGGO4InoklPdM+ArShSVgdiMij
++v/Eg8ilwI3T4rNjhLkBr6tcjZBU35lBiZVNhFlOwgLAgUZHyJ5tuStvH2bVQAPeIvIErZwpQlf
b9nMr4FydIFLO9VB+Yd3lJ6lgZ1jafU6IDTsriZ7ISchaSwAWVi85ZM24T2ERFCQQXnnhl2bPsnv
jAHhQLinlaajW0ww7dEnBt4L4av9yel4xI1eWEPKlqT9dQTM0OXVgQa2a/O1/hp2LzE9HZheGu6p
PbqB15YrZIFnSCqAN3Yueruzvt7UGqXdro3/EoURuuEaMsOOWqfK3DEZ5J3jPT8fkNdD2VbxRZLN
S4SdtdTu4RRRV2NJJaNqTPpCHsuknmvA2f+iuirMVCWBwJ5rVmDBMLzuw+3heo9O1bakqCJg5Xth
pZ1xku/4vP9Nb0s9j35QMLGUnS5WqkGmcXf/5OPI4ssBE+isZytpSP/bk9zsvSuoVsXsV7uix/ba
GtgQzPV2CsfZMtGqNFZ4A49h76ROd5mp0LH3kxfONmjpf9Q2zLPQzYtf/H4tdnq8OYYYVGlEUP2w
Icb6Fk1rHUPxstS/Abw//rui24OObcUraSoxEkINIxj7EReo1hJ2YTfZl75Hm+qQT5kRumpCFyeh
6GEc45VJaLD5ev1NqlPzHRusumYQzZaM3LW9B3mq9yCHbCsVikWUEw84piyQZZangqqcr006/7Tw
ZJ9N5xhNXrX7zkXNK15LIPP2lDM/hQO55wveEBvIYAH0VM8NLuUWuybM78Hsk20qsECpp4zGX7nV
E7fM4IMHnFtNL5G++kiHP4JWschRvRa0tjvTII0XOlD1WeUZ/HX2MLjC6rh63HS9jrXTjfmXvS4+
K5S09rCI38CaIcTDvLj/ounk1DCbpsuaAFSkSMdXdPbwhVlieBGts+sbyTv0rHz1IQmsmbbITLAt
t30H93RvV67Z0Yk16a0HVZaM7iFtvTCyvLl+vCyU4nBBwljVAcZUipjoxoRW6ebKczTn6tU2CVgN
TAETJPgx/dCwe1QBY20SbO+Q8kndWEHuidvXvy860VFjBJqWNX18oyFSiz1u75fguU8q63qtwQAV
JuGzHHx5lqzNNqppnj72E59tqRJGvPsMw8U36Iv+ED46b+p+6d0D5+EAK3+v/pC1tiISCsfbWbPR
xRC5ud/7d5a7GRYSAvEc/Yf0wayTm24GZ63axkNC/6rDQSg98WN/oBJ0IgFXy1lxVcMlrSL1oAPw
2etP1cjaw6KNVfoLhYnvbAtBr/+7uKppABOMUExgTjAtzhRATABXKCdQwZ2UwixJFCR05vJ4K48L
y+vmk5whlT8OnfA2Fl5ng9Ogs1vZZDCkC9YemIIWeu8mZ224urNIJSfJ6NGyb2dd9zN4diLI1I+a
zaTgDg8QxZ7HbYTWww4Pbd+Uz4B6QDM8FT/+SEw6D34FkzgV4TKLwtXiDLICU3UDfxgTB2tCSrkg
Cn9T4UNDGX4n49pH027IKy0l41YzOWw36bH0OAQzswYa9Lfy//e5Jo/Hu30pK04LWbnpchVxDv59
1xDGRToKKLY4eVfygaYFJCmQGuiNP2zqssdXcITPSD4GHghDyMWj/2ljnHqPN7dnUqqgd9aXKqNq
BUmg8PWw8HuLWWAump79YCytka0DES0Z1ldl2kCIWKkz+RXXKbkfTiKJ37L+XKRpE4PbofS0rVpG
21DxdfXX35P+8BLm2r8DDGsATuW+VlYLLIS7onjmGLLmdzlL/kayoF/GaeQMmaYSvPu39Nw1AIvP
Ku7vuKbHsQ1OJEixjk6mQMSLX3G1D8ElB/5GMSU2DMwGMNpqgT4MFvMr4AzB3nIKEvnKtmIv3tPh
MJhRlwEraGTlX0snclfezCvptHXoGmUZ7ETWu+1mod85Bg6rUsYtfVoE6nzPW/c6goV8oYB4ZIuX
EWYSESZDHJ65bruHnd8txUS9Bi2Yr65A9bE4Jg62pDeCRhQ9wLJDDdxYLZakAx2v41WZOCGmkpMj
WP1gSxrkfJbDnkLG3JUvir2XaNZVQiHtoJAvTMAMqEbonpFjUUqrIO8jtmqKEhRE39daPRa7pyMh
bTlOE2K74kzTlroK6lRM3EM3oJBGOlpVCnthRZmyDfvm8FZoZ91qVJLYLG0DOOE/xg3pWuKEZU0D
eS4gHfjfZm3z/ei6bRpyPW1na0haCI5+apInBNBRe6Wry7CzbHiQhQdr04KsOehj+J976wSFgqoD
ifZbE16W4gVdW7pN0Hz8lSaUTuwybMKvxdyzgcRojpe+tlsaO+jMZOWqa2rm3eGH0NqZOLhjkcbP
r9wDxnWz9Y1jDEZCHbZ0Kmd8Wl5tICQ795RHmLjp7vPtuVoA2Yd3H0f9EuYlCBG4FuPtHKh2a7hw
RvX9h4XI+aHpQaePxBxpdMpyApQbYgcg9YV4rb5tJgl0gzEwfy4UYU0VsbHYFrpeGkP0C6ljmwKY
Rha3EABKcO0Cm84yFf/ce5MtgV9voLIriiQWrWOih69IsC1YEQ3Q4aajnhjtxqZup7z7vcppqsPm
96MKI88dK66RYwm5uXEsnEliY8eTjhtAYaaez6lh9YNyD+0psufUc6zNBOuHf62uPFzxppxZDfy+
iqg1dXfziQjhE/pA0uwDlZgSheDffZ3P2N41MwlrCwbquPM0ARJuK+IyBJPHosXvqirRxBu+tKUM
jIv6/gvkcar/lAqjVReYLZAHkexSQDP0vfsmmO2D+BKbq/BZ8ArdOs34tjDlJsW7eaaD9tRDFwOm
vRAoCgJg41pt0EfLDK7khAzvClQPC4VSrs1MoYaiAakA8PakuCaKkOU+gQ8CU5B76XBwaYnsJg7l
k5oWm3v6zirha5l3bta1dQUi6HYhXMGVZyV1V5l0f3EoY7yqG1yHKXoRVX2zNUvqR0qpIQVb48VG
uJG839ci8/0+wmXF5/bY2MWXQZJXZ1jRJ0HOoThH3CIyYSxDgcU4L7CK/sSbnyjT00g720Zvq9J4
cQjyLOycUM597Vl1OUPdPun/SbsbWBDG3PG6Gz8TjS4zrI4Tt1OsajB1ekMYHbs9kvUjOItT3xAL
af1l6xaYYBHwm49DRSXpkwSQtX5drgBIRZjHnHOBnTZNYRHFTZOaeBnWrdKjF2b0OEf3YjgASidz
jZ0o+ZuMqrFpyTdQw+ORF9cqKOnA9rIzwnG/cYXs46lOMfPfRnc1yGTk9/MJe5itC36vZ9XKhESm
ybqHVSctSlXiOPYtCxUVe1Twn3EgK+z0fpy8cw4VONsm5m1Hd2s1yVqL3GFy4rvy4u/oIU3R60+n
xErNBLPVbaN4w8l+xwapV70PHcJM5iIIPi7bUiHyOx3190WW2oaM1Z0rSGa4vNoPgaDXNAMof+RG
l0AUikUml88Y7I8dPv/52malD9UTEa3pMt7Yq/83iL/sAfYmBKzaedz5sbFJiEDBJYNKbfMYkKWh
oDe+zkRlmuFz/0plTIAb5uO7wh3ZcpMzl9q1sLX4aEi6Wrllk3I3Iiv9+G44+KDItAzWVJ/4ZZJ0
2GzzDmXlAm5LvWXiCvdqFN/8M2Z6pAoU2e+AEEGo8cTNs7bGDAc3qmN63zVHCItVegcz8NfqsoxH
VN67W+auejJo4gMvhGF57owGF4GHa+EGL05LaEKUQ6ZXGF7NC4NOpzq3oM1DgGHPW013yh8fgc3k
ZaJO9QDhT5ZM4pegqJPZgLa+M8xgydFMjRQyxweXnoTjRyQFAcNtQFcjGk8xVixRf5DoW3hnRI9X
af6l2qUon06rjeERmhyYYIYmRnc3ylz09JGCdswtxpgDyKm+JzvLFgw70AP0HP+uSDAK0r4MGlRJ
3IJQ6BZCz9SpEBpvHcx7DxWq1cuVTYwHafzcbxR2xBVlZxBQyH9JSp2f4tOSZkkLFe2bF3hhkeZP
/yEBXzLmswXcrTN5DXVcAdlBdThZT/tbmUA6f7PpKfIKNo8CNnak7EF4VwMzsfiH+NBxqIYZgIEG
GpLG9aBwj0jD8yXTO2M4F1GXNDaLNd+rCG2eBO+RMZFM8tfj28qi9JEBkM5UySF+n9eB6WAFvoEF
Rh2ItARC1tsBHrFKfWNM3hemQt8ouBlpyXx66ZcJWa2uUvr/VQm21aXMZGAXUMSr2N7sqr0+x469
JmLKo1oZsfmM8dtXIu0U7tqWjY64mpmTWni5OobvtNkPE1Z9O5Q3iu5uDBVhshgYp1fw94IV8Bly
M3vAKiHKyUaLhbIt8iZe2B6vmU2g08/t8wZZEhffZGqOvhAb5ObXoBTnpTC7CZIItzbEf/gbicqR
Yx88RtO0vcM/D00ATOWeuEWXt+i+iwtEicdxYyQnrsOmu6y6dzuYNjdOVA82Eb+605djY4ZMTKqQ
qWhQdM5+oSoujCCw1khvITpFB5vvRY4w/6qeKwOUzHxQh9PvjH/SZggPvrbd0Peh0sm5kc47RBS+
9L+Geja9N6Wfu7MMhVbWHV1eFvwiMZl600KnszUu3+MmMDBzz7dZzC/naydXMZot0DA9Mnxrfjsz
o9rx6QvQBGRudN3KnEWMFtkuCkp63Zuor1fw643NGFxjGVTOfxnGDm1NwlAgT902tIkPpxnTvJJ3
ByNJwRcZ4t9J9KsUCpWdPN0I43ibAdexuMmvgbtvHc85UvIBzbvIKJHpxfR+0OM6Sy8cUwmjMy9d
eyUbXlSZwHr/ZC6ebpfPuuvq4xXy9iW8ymNtMJaPTIZQ1yQqOoj0jotDPbyVEhaJkpC76eQjxUPg
p+itpLqFUvq4kFyxDp0L9B5RFAPA4PKYMbrleUgjEjziMA9rnGychiGwigmeB0A+wFzaKH5Gb9xs
YlI8m6NqxYufo6w6CmgtT4pu3/g2r6WlBLA1oXakg96VKIqvUMM5I3MZLpzsrypDffGaSMwIBiBM
rD1GT2TQFFZIJvZDEjLuuhpIJuNCGakAL5LVI4Oc2CWFQiZHVe/Kl6YG3DjaPgnprn0LxR2I21Y2
tXDoz8o1f9LuPZ2zmCfSa+6MEHcznXsuxlBX6Xf0XamT6mZckAWwZF4DM/3QCVbh2SaYsb6mdGl2
ZeY+RfN5i1KxT1eKoWoazZfvfmsRWkWN64aYnuPn7yExC5wBIt1kAYDNqrp5y1QxPS4RfEPTNYyV
CSBGbRg+ZNTyplZR//KfnEsnzSjn9/OAHWdMIPbyY5/TWdk2dhnH5KCWAwzkOfhu3oHRoygOKIrA
qAgcmZZgBKTAmKvOo2KLJ0AkJw4S8LZFkpRPR9DMD5CxkbcEwmwCGujkVK2AioQK9dWj0CSlZ3jD
kfg8vsFlTUgUvogSnnh2LfR6955sOoduNfZ1li/dznEQA0wyikt2UaExp7IWEpGEz+/Jiepz5jeQ
PggvqHLmBcOTKReyU6EfKsC8Dpir8a2sbVZdrB3nRoL5MOK6oYfv+1gWr9bEngJlNJ/CudiCzJWC
7nFGuvN9nioXmpVvZgLtbVXeirWe5acuYWk0G2Wp1bODcsTHv1QMbsov43joDrDqpBmix0OaVWnV
hWNUTfXd2cyD4QOGY/QBRcSKRUDEFKyjWmyGr+O8ICrk1T+cOzXTZen/ftrlWBsMPfQMw4wtVkNV
7KdNEN5soKluW9VCrApPz3p0wKocs2BkoKmn884P5eOJXtaz4FzK9ssAs9BsFPEmZ/VR41n5TVU6
bu9+qcNjWCqm+ZYZzfBN3hNJTLe06MGyP5RAMYZH37fzZp4qKKOUYY3HGI7bLAX/Q8wc0anFDZPX
Lz6zXfl+0X9xp5kmXycKFc8Yq5w1Po4/88pL3GfaDjxmgZsIxytCwVWlIDjZlJMjWr6hyoQG/466
1Xxm51sQbmJWyjEamBDH5JZf3gFRJSE4JLNgeD6MVSrOGaB9QIwYztz6HVpmMRFKX44f8rKV8xRZ
96XmM8m8ZW0HzYgxzwb7K0oE7VkHMzJiX6I4whmPCk/wEdahlv5hnEw4YeOqgRjPzN9LDSXPZLxR
DIUbCD5olCM9WtXJrzAw2Y7e4vo7P5XpDNnj/c4dR+OiQxzFj6XaxaSXnqGJU2MJwo5j9VLJnt0W
dUoBH9lLiAS1wvUh1HpMHiUo8RCmC99tAupOvA2dQxIgyl5LLT1CAD7HH4fPH7Cb6jJn9hUgazAU
87/Gz0ukg5OCekdnTB8kz6LlMHv2UNrXeCHpADa634HlSOgGXq8OpUcxc8f6WZgl75gF4+tLeSZf
hVQlDN1KQPDYwUCnE1TWEE7oy4ieJ65mJGzEl7tbzYQc/f4/eU6xGvWne9hQM3UjvkxPv+HDpjqk
rEU8PuXSrU6DlqPyUsh0H05odlTQEVl6x2rYLSoTQCdSHpj6gXxG9VsDBbaAHCEN5cMr5aRwds9i
Xbvb+Su9JBikr/O9VDQXGZYQE4MFeaEANglDTqyZBkPFNUuzlEPF1XnwAfCPLcdjZ9ssDzZ9p+Gy
vnHFTJWf8Ebq2jTXxhPmRjBkL7I20KS8CHek1C9MrpGDvgHrVoGeE8QQmYxchHabBvykerXOLJTQ
A+9vyyVpCR6AXM2G7g7S+puTVKf+RAmaudrH5RKfLJCKcPoWQynyd9qsRJcKrGx1tB8flcKpQLWR
8J9fn8pW4aQ7WJ/zel7KTpZhsEi/qHLBKSTICH3t4l0I5pft+Y2dVGVDekNYTrmltyFjL3obkcSj
zCrKmM5a4rzJfruxWbIYQb42dtt5wrxbP+pxE1S5ThJGBLjNb3tk0sF3rbcm39FoY2CQBifDFvxV
r3ibp1N3k2D3CxbqfkSpYUjHCNaOb5KyNvBpwD3Rqe71SEi/cFjylS3qPVq/Tp64H+4eUlraOdvO
7ZlSB/p13fnPEhXTQssHI5SskzTjogtjSa9hAi9qZ4MBeeS+OoKgNpztb2eIISBQ3p6WCX5S4W5O
Cn+EvqARGJfj8DZ4zMyKx5yQcvPMemTUpmt7sPxOjUuh6aaecsx49MqRQJ+S/QGwj0g8ghWFKHi4
fa4WCSO3vWHgIaSqlSFvDIKq6nhIo114yMy92z11HwiXI5EUA/nP+GzS9vuf9KBuF7pr2Yo7rxob
BeITKi6H08uuMhp+f5c873jwg+FuqjvzNPEOlEDWnCpPTbt7e29Hkwp+aZ+7UMZcIvnxLMenVKyr
apwBbM0rRdG1hEGwyFMjgA18CuMQoRRA7ncMaLNZrB4LE0dZupjBe27KEq0qZPRPVn0QHoJc/vSl
GxMljsDPE8BQgJX28efb1zwxWRmWJbr6GOw5m1m2uet7XohlnxfAtvz9TceCbl/uBujIb4o1dvkg
ZFX+dHjKksOSU6WrXM95yi5N7LM0XSUAF+uczVedkYuR70uDJCqu6aYFQX+Wwrlv68HCbQ78SCcY
qZJdscDgO0Eivx4Mg2/CQrBAoNSqiQs80vRaJkDqxaeBpvNu0uCgFpqXzJyvSDMaSUnn61ueE4og
hzb6GXOZJ0yOlCh4QOvBCRpJJrrBCaDnpkJq1qfHlAkm/joWronjXtsTgary/qR1JUETUtp6J9uY
oCfQjHJETZIdkoNnL4thFLBWF/Upo3iORpzjzZ3HlrYLpSpkliDAUafbfg9O5nykZ2n8bRAiINA4
A7hrTdREO+KSYfRj0IuOhc1AYlI7611cq6F+flwM43H7GJJgOiEde2mQi7aoz31QjkgeSkta3e3v
b1HksuMlzyUXUSjy/9s///uMJ/ycJQ4hN+2XR5+8hkLB75p6sY1nuzAjL9lbQmIMeUatYxMIN1AT
nO9Uu2/EnC9bpcN7c95oDBd52GSnGcoeFGhcH5wRjx27PnXlpi4zBnV9caR3UuNJJQNv4sgadERs
jbfB4Pt17Mrk/0OxfZd3SQJzpZeROrRiPDbcRdMnZDm2gb7LTwSy9SnKb0kWh6dHHTykDiDfRHrw
PL3++0Alv39cmtHPG8hgSLrZXl6pyVILTvMqWhP8umUzS4Uw8QoqsLmFCGLsR8/teEhdeymM0Bpv
kLABRqABTaWYS0yMOOVaLjWr/NtLG+rdHKjWM+gb/KhEDhsUm5vX8hvN0DAU5ef272vdbX+6WNrd
ClvD2wDAH9HLV+w0izwryc9W5z5PfYJRJ8uawnoB5phDNFyqEfQiOsdLA2JpT1NfHMk2gNisJAYb
mAGDsAwPC+2KIUH84Ubw/yAFl4o92fo8W+6nJ9NQfKX7W4cbWJk8XEJGv55zgVe9Cpw1Y7TtnVgU
qGRwYiySE3nkNE5lRV6wBrclgop97KDmN6UPgQxLKwf840HcoG2ImNBUPURe9P9DE2tmWBhQg9X/
fJAlH7kwhvy4PHiz9VmbfmpnM5P157tj0SUq3DK5Oz58rCsyCrPKdhMGcLfY3L6SANwYZSWk/y5W
bb4pb/diQwQ5V8CFHtC32J9SvoFaFCC4/gN4wrWWH7yTcuXZhkXEQEtO55PzsdeVmi6zSjh2vXFX
g+2E/+1viXhpVsnRtDXkIGW+/Inzo9q9dCe1OaVsjP0OW1xxGinh+zYoT4qJlS0vt3ArT185GNh5
9jE8ty1KGPPBgCJvKAsW2NKJp5fjQu7a2xLf04/rZZmG00iDRrwjPO1rnfgnAfetJvO8koHGaplC
NSOQ9g9fHfDqBF0XD2SywQHjM1Ify9HnlUXsweEDF7DPZa6YAy8fcLeLwfZz2E2lKIS4zrXPRFBz
QNA3nEevWj8Owg9UiK2OKe6PTb2vpDGZdNI0BU1XJzgvxkfWgSRx/D9LrC6W0D+pNXhtVLF1ImIt
WFXfdSeFCDtb3oTeSjvCywFZsgZdcYdvUMVLBO5YWb92apzjXLwbMk9SSDlt7RBxdShZ324f3G8i
RId+Fp5h6uS/l25pIWH8er66+JQ9S8hSVd8O+r/3XEakTSFXmauWIBGJAUz83c3mZy4Bo86dVIhC
Lpxcdy9YACfmwk2drsA3+kIdUTJ+SzFbDXWBNJL3YYR6ogEcj3NRAPNm6Fyjn3dEficD8Ee5hVhh
uPjpruAvoKKq2DvKAVDrIVzer4N30GtBsTEYa+ygjkheYkifbVcbK/OSzbL9jrKsTc2rPhNyi4bH
gkItZNnJlxc5TS06cJ3pdpu0yN7ON2N3c2EgICBsxWyrRt+w3eczpQ9FHRrAPTo9eocND44yJLLN
95HAZ8KrOwKw39ujVQaA2foBs/8yCKtnG71BdjbQIWOXAUtzvVfKhkIxzgRr+Nvie4nrgKCNYYke
XlC10X4noqH5BdxHJRdtn9r/a450khjj48RfvvMH14dlXiBbT4Fb5AvXe9HtCAz8jku8NZgss4HV
skmENSqX4CUjjNd8/SFjM4KSRXF7R8I5rwbMvBrRgKX0iRGlrGCwi9c4Af0qSneAYDvffwNHV6bi
x7soW1j3GhQpOxD8q+/YoVLraYonAA6HoXV6IsEEdHbFCtQIL149GVCJyQFaU0Cf44Z1Eemu0APp
3wWTxut03pMOt4W55Kfs6KdF2a8IHq8XUY8Un+1xi4G0JSeefUJItmwYWQEsR4DF4qx1OP8EvFU6
u1hZK9Db8IXLe+Aq18cr1lM14WV8/rdxGYuyFYbdYoT9xigHOEtnDWT9kHuml5JVHR6zlrm8gC7E
4k7bs1JE7s8ctOKGL4eO/M6EA/AqbeBG1/4Fnf+N/iCf6LLyfZqvNTGjaRrzATBTgkPAVWNkY9Sy
TXpkgAP+0hDfMs11G46patQkUGre42FWuVlq5T1H7kIWCPcZB7U5VUtbLcs3a4J7d+lvn6GIJMhZ
KLN8IX8DS7VetsMEwXyt1c8xDEv6XajoFAanlxNiyXGTFwFMjbcJRg1n0d7qT3XNgCALVfNdsDT4
7/xLPVgshXdOykELktCn/vqHy6y3IOLYr95D+jqS4jX2V6XHoEj39GtWOiqaeoZHfCAXvFyQbFnS
VSOvlg4G3oAyxE/ypoh4EZRQqxf/qQEuTftyihHtxgvRCoCPd16xF/9dn7ST24MUMruDi7jMy/2F
ndbbLhXS575rGHCcYiK+hxFUjKwJqkR3iJLKg5lSTyUyCifvFfXPDsLVKDGF5dPTedYsJXhC/1m/
L+bPfV4l3+tRLqAsTOfFC4AAEW5901wzXmZ+fNjHPgTkwsK9X2HmBhWg7NhAQPeeTlmR/PUxuWkI
bZ2nIhwoVgrFjWihmHgyFuIjtBjEXZqhfTYZlRpzAxQPN4Iet0mzY29uesvQ4a0yoGcsIEoDgnUN
TRsqbQVnWOx/aA7iEwH3lG9idt79QYxfpg8BrtNovjMjBHLT0ij9zwBNpOBPtzrpseFcaB7aq18w
TArQ/ZD6zWBHyhkawypV817ulXr3R6k4WGJ24SKtJcIwE1e2NPclaB6PwALyTqAbioz21xrxYc2K
AXJb9lupULkVdqXk/MBC931Ht0ywYX0MgpfYqx5e6wm6lFXfy4bm+z5XgOwJkCM4Quq8qcmVSGG+
G9lB4PMTrUhWkh9xIlPobYdI0xbwfTJ1RHX+0n8QeGF9XJwlp3Ba/EoqYH1ZHBXvrXJt7BBkywmI
FBKerzsUtZQ3TKrFeiGk/8S72rhcpghoeWqxxYTgAyYVMiccvuhsZycbUG3imjgD4SwAwC51bhYC
vx19NynWiInpQagazo2J51xLTsqGPZ+kkFzwNX9EN0tEZpT1ga8LXt5kxLtNf9hIMf9Q8WSNVo2p
KafcFdEsl4SvWyrOza/oxNQeBGprqMbxG04kNaPqMMnO2Fj+JEx3ZJI/qfwAmXh29sAfjxXatsuw
vTxR2Ji4TLWZTDR/N036YXa+hBFMZ0YLRlGa7jA7fvO3k1AIE4YWK/TV9t3eZ/Q1IEeonOKeURTb
PzRlcftoBlTBWX1KwKtk1rr+GLzvKLHh9ut3Tg9m/GMAM/Ah3kzpAF8znQF59NtxxMWxJCACWogs
7ZoT1ZEX0Ehx6hYzZ93boTWNjEn0otvJ/2dzzU8o5FjqtLUl7rL8vqrT+Jrr4aS15Z+Jg1zyQ/LE
H43HTUGTGRb0BuB9OTrW6hAIWRptMMhpyNcCvYuhdjjbvaGliHsDO+gGbnaz3G5bbJ343tsFz3uJ
M7+PXdw4AMCEsRHS21JJdMoKVRF8i2n4mQzGOZEFzJ5SQIEL1MsRQ1YGpr0rhG7WLpRDhnqCCwfM
OCgz+5xkDpM9MwcJxvSyD9cTATb2QRHdE2j/uxus/7RLUBXCi253upYFhvdRdlEjrAOtc3rz4Ucj
zuVxYMB7JU4JzTPlX0NC8FMT+cSLfM4fdZhjOySuLVAN2M27K/P02kS2tr/cC0O7FIf/aw9deLxr
yoDkIo8whgbpqVeiOlCYrtPpTi9JLCPv0mxrzuCJZIDJdY9iHaiWzZxHmjbL2eCyJPhfwXPl/Mqk
SejIkZJeh1dy/Z0gKCnAnO0yExfCTQ4agXgNgETmU1Sc7dniHcII949wRTpOpqHiSzzEjgaPqZZD
bHNq6ST5DtsdGQycHvPajv6oUv1TmS4m+tbOopOz3fvF9QPbf+9xewasR8yoPOdVLCjiqi5YtrHN
jHtZArckk4kNRdMWw+toP3g4OtCbETbZdSAmDNNTWKk3qtugIwwNAzezUTPw+4/7dmO/gQRxggRz
y1+/IyChClMRDVBKV6+l41guNbXWy1fAUiKxxGIBisDyU6aOsVUSSOGKVsy1E9B9OTaruR4Q2Xw9
6BDjGxAejct5agayCdJAQAigneVzapR1rt6giKMuu0+NJ2j8ze7zYML58/9s+MmkPYe4OHpPvqsS
/b8Q5+9eoSp9kwv27YjMZKYMkQFShLT/63auGbUE+D7XUxzkh6/2DJJHqc1BwL3nnLrigAsTDalB
LwHdty8qG0nycTeXnZZmoc7wchpaIhRVevFZPq8InqzQKDo2uCzKf03kAieGPFD4zsF55UUYHL1q
QwvnJn0Y+sdhUnDP4PcQc1onKW1qiPAS3A7qODlqCxXM+yjxwK0IxHZT71kQroSvUMcugkb8Y22V
2DAI8PYMXzPkwSegfk5vXtiGio8K3TO9SnXoJ7mI/Kt94dDGzLwDXbbxXYHiVLTUr4t9Q/m0mgKa
WrvzGEEULOsygAjupSeYScfMlWjb7BzvjinaOCh/lwYu5R68BHbTUHo9hvy9gxNoqUnSSEpX2k0D
o/6QgwIeU6BXAwscD3Jhsw0fgOd8U8w7GIgTrRYxQIJeQnfZJjmCSvtEiixFw/qa/trdU5qRl3H9
uXKg+sOWy7p5iw9p+so57uSUJjhHYnjmu/ELBWUSjgbZJujX5hUIi06YS+I9M4rq7SaiEE7M+rUu
KS0A/X3hTB15LXZmKHLFPMXktG3B7nAItTbXki4B6q4/C5XXMgF4cOolmCwRCKFgoRypJNLZQ66O
p8rDOcuZZr1UbF8nb7iLD1+GK6657dK6Y+mXRUjOWO1NVfHvYgj/WY1P8vPP3DdAUvYKjJpQsY6c
j6TeNdjCtS5KdZ70jYgB3KP/4bY/BxvKE5gX7anhiIfMQUHypk9vF7ifvGk8bHwLq96GAwa1/f88
uyIcxEY9MooNsU/Ic7RyQe2H09XZBD8h/sQGLCDI0xt9iCHU858rSxFkWfVCievkOxkXMuvxgJlf
zltV6D802bc6rij2kgWLigxFEbpEsgP8qdvWET19gERaGYP8tR0h/fzS6mqzbdEA5b8eGAKaJEXP
Xm6YniSwB2u2GvsdLbPTopBlCWjOQiGRhR5KwhYEYoOKY57+n5oYz9GFoX3BWPo8OQuU9D105KGC
/YbpqNFR0d07Xq4h1LT+Is3cfI34NfPZZJyx1KZavZcMeaZXzmAysXQ5ke2xoN7hL4z/bmwIv4Vs
Ee/Ad4A2CP0C2Pn9+XJFyzT1wJTAW+tymBstxAvbZrkQfU+aHtDHpEfmHnqEXZYKqnciMlj3IjP8
M7CxMjHEENJCPjeugyzjhARiSNsSj8vPip4+IPVlixoVASKPT5pKustE38xLu33PlunQJDbQqQoq
6+vFbYLWjyuLFDaela6b45FHDuOttOlPF6873QkJkBqSeSMnCYrtfz57LN4MVwXTaPfASR+7kMj0
p/904cp9vbc/x22SpOn4yFMCnWw5IF80LywoyLpXF890f/v+0/y7tk84xb8lF7LgCz3uRqkg/6tM
N36H4JzSLoKX1Qnue3AoZaVjNE+J+z2jNKxzwMYbZdgyUvGellmhAkuRXnzL0h2yr8NE4jpFuk2W
pwE+BaCcSbmJ7HwcmuqMaa9QjHWBs6W/tAzyu1iNmatSoWUQJnPvij5JiUBHIsxFw5jjcC1Qva7y
HNBHatZmxGJyI8CQd8empxli0+4pinb1qkEnVfFk0ZlKJ3imEVufAtaWsN4/UqqrA0uPWe1odCjC
udCf2Of2UdBDQx8KoAU8hyz1887hVykG7/O+pBhgM4ZBi8IK4QEDo4YH3BEKIik5eZ02cPgqqU9y
f6Svcp97iMmxJKxtZ7yX65WkDPn9lKSx2A3UZTUPFhPR5hN/Knl9WDr9pI3E118Ww/tqJXUgK7p1
AWSgXeIjEFdSuT1DGsNZ1XBVvYXGpEIvT/AN47Ln3FlcrsgDmneRHT/lyJcpf5lgGNzCGz/WxG80
FkjuGm7CBHtertEcDrD0Wj8oCgFbmNU877WlUEGaYCGQJXOM7SAL3bevFUxsU46jeU+XyIq+CVY6
rX47ceCBh+uPawMZmrqmdznG7h5/8mLUQS1J3ErIYakO5cFMhsbPn7zlvabGYPBLPVYizPuRE7Sq
Qj+jJKqYMPmkF7GgUaUTSX+4bbP/p2rgZyp7xWpYSgWtXgDVzXsvfSv49jlTOutIIXmLPZo4OsEQ
JawCI8DvP6H0MqKFFas2P2e4ZxLAjwM4La3vyN0XQphaWDyUs8he3KmCer8U1VsOUqwioCmWFV9e
xAQ9LT6KFf7GgDv1+dVGC0OiO5lMpc5nNRhmlKVjxN2Jg/PFuT51wQuMdLZkBpBEHxR2mPqD6NMm
j8pVZGU4Ox/Y2j0C5bJwM01SLI3Xl4J9diW/NexOXlmL7mAD+0ed3r3hYSS+ZvPgUol24mZHEc7U
eGPat9ZHTffu2H3NjYgl7br1zLnNYgkv01zB3l71TlN7nOTfXgZsALFa5RSxKXFW4ysnquYh0yS7
V5nkTyTWLkuTaN8KbqhHCItZVii19h/Au0Yc6LeoEV6bY1908mm/V0iUzN918UW/wruz0l3EOl1y
ACJ82GP5kORY1Aka2vnVyn3PFZiEA88Ui/qS+SK3Z7djI2oFlbI090KU5gkqa+V9YbZAiyuOS22f
N1qzHeQW3/P4pNIFLAZ+lFQOQUACOBd7UG0SnL3qbcm/9sbQCSR5EM9P6nY36ExHS6hnG2JIfJGQ
Vru6JihRjbSM5qvAIJj1qfwMqLIC1YDhcPA5QsBQBVF+Pp0Qu7Pv2Ta5TxLTb7WLeL0PeK/x72/c
31nrpRU4uSkkUpq04OjZnarq/T73Cyexa4KHaKsllfyeScK9tG1654oeEoo6GhVKMzJhtm1TBHMg
7jUQIxadwNComo1Lb6fDQwApu0ezu/ls6KDHBjufpchUCbaUxwAr72Qv25fR4ypEDigMbIF5Bp56
GCWIwbW/3ik1ZCooIxGaqh8S6zue+KN0o/Kwrvu8g18Tn00TsmgPyZIyzpSqmVoRJivEN4ihKw2s
aYqLn5yd5HI7bmq94lag0gctUugFTG4RMb0cTKYMkbwN/maLjo9wC0/Yum/tlSofa4bwHKHjdgFP
X2itJotYk0/GXGl7H1jxiCAQZd88Npp2rtR9e6EM/ToGTzGGUqy4Q0lVtT6juAypKQZ23jrkmcXg
c4kT2rl54np6Uvry/BWCn0uKgXK0kWMQIdx6n6UTtCdyqjB36U1KY/eDY7cHvFQUCtTfGBDdQUJS
3/PiqIbfl5O4QkjUqTw1gS8R2wDoLjG4QYGU4Qx7oq3bJKwmKMwqp/CICImq5ufCJhT7YjkRfjIJ
WH2duxrWmrD9oesHlNee5Wjv/LiNW78yQ2ImqUeJIn3m4pcqhGcNB1P9WHF5+OnJKxFu8Q/BbTO3
ltZeSTR3gZcIjhICh79OITNPjaci0Hp0TYBjBXc62Dg7ktgCcBEQmaY9KyYWM01EbmJGfLjYjUle
z4Gp7kXQ4QT5FKDqQj+YKQk2hXIdGomHhtdv3GFIz5G0XUW79mIw+++iWxYlTSu6AY1HYZV5yUHW
wYPUxSOaq+8jJ0213PraMJXMDCsPhYd/jml9Ekpxam/iY2VBD/I9rFjfCvNxjzu+INtaej3a+Usu
v5zwIkZ+EhvhJuClx8uDBhBMzSDi0fEWp/Bg9dVbhnaFG111v8HuLXetE3LqYER/kntWAgNiVprg
VvnNFAB7aIIuAQgf/UC9dIVCowYnNexibslOzccAH5/0M+TEbgitoirKcK6x8FzC5lKXEMivKmlS
msrZN7Yf/CxAkjzvyYY/TKvDtU7IF3/ShKNkIqJCFuWgZwMZE/gBzYw9kp7aZfa1zI2OFpeqvUNC
LSw5QyE0BtH+L+lp3I4agCd5rTJh/uDmIG7xsdMaUpmmyrFb6QLXZv4EPb3nenROWj6teW7VGogG
WH1rmjYQBuIO6o+Hd0rlqcfU5v5XXBBs2diUga2ZaOem0ChDN8gIsYlmMYOd/f6mx2Nnor8YXSym
TWk5D6OWi57RNJR8dsCVmzl7ZRpJCcagXvmkDfBhA5MyfJKBk/6H12m+7jnM950BKYGRhMjp+xhU
z586diNOkJ5uwkJT2mHRNF8DtX+mHGzFdYuvOsBfKom83WOw0Alyj5RQQO15ryfrq1xAuFS/dmNh
pYRrFENQbGuIMHyVgVuJoNMapi0sj0uXYh2jml3vJCKt5cs59PJaflwG2QKrUv9u2HNAkhRbwpo/
y5tBYat8K3nX3N6qF9VpudQV7v7213JJp/NfP8sFromuzfPqxPjDj8ZWAGXkIz6EC4Sy4nrPTA0o
/PqgrxtaVF7Ie4E3JwvL7XOh//GIq9o+cjTcpz5m2JYE2sn+rRXDEYie8lRyyKyy016YdbL+oVRg
GqiDburNhYDIr0a8NdCJV4hcRZqLTxWCGlOJpWC9Di0Xffe/jiLYt04UwTeR3tAXryaGwJe+9QFV
9P2W5R3mr+fu/bOgwAY6zQLxRKff/YUzuCeE9mIYuewuRQp70CLA746LTwubmjz9kwk7bkwTgT/x
tSsJ2tkmN8AiZ3drG2MWIV8DJtJ0XEc/Uz3U3GFoVq3B9M1f8fM1pF60d8InXgqC00bi71ULnyu7
bGsXVeDFrTOdXs5pm3tRRscBkABF15osSQmli318eAME/E+8ZuJnc1jAcoGWqtVax0kTenLT3kbf
JOprDC2fMYVQEx0xFUU0XErDtKfSV8gb2fWeDr96m0oqVTxDrovv+GPFYWeprxO6J+i2LDCvuc9t
5hf7Vn5kMUYNJn07+uL/W8ulWqdCgEyHlFVZ+6r1ZdKWhuP43gu2OE9dTp7spV6d8ib3sitfC7Ry
G7zcisdshGypLSpzClXDUjxjiviMpQ28j/qBfX4Cwiwmm2PIJWKH0Hp+BeHF06FkYy3oQpoU2247
qUGpoDV94rT2IRW/U8oyo+b317XdeE1/4W6SiWlNXDskzuEUEdMtsU4Tu7HfFQdydn17sjkEo6jI
7eq73PlF3nJDNpHY6G4J413arVYG+reQVnm7Y+9hnX3SNg8K+x/SV9PlvKsj3YG/2elQE4GNXg8r
jRyPrglUUgbxAMqPP6IbNgfs15RwhkWmNwyQ31NXuZ3M6/5Hl/40YTC6MYlgaNisb3gca+QnxkHg
T/OXrOhWkc7Mv5LPqomhEhBoOFI4b8Fny94N3+EXmbXZgsFYaHH5d6GbZKpuzXRNaL8bW3izQncV
8OBxUhZBjih24oPX74ZzpernXZ7ibGDYB6aOK1G56x20FzSCgoipDSZuTdanLd3wJZEnKCbsDJlh
83dnvySEC6Pj6SeeWCIJXtyK4Px7tfyalrH9pr990nd60p4nijJ2JcvguaP49hDl2FZ1lm9ajDCP
9z5LEPyURUDA1MmdgKxJSJvhScxz3+V9r7uGT1cvhiH5m6kHfM8hO3iyCEXWe5hbGrKAcit54rFd
yAOz9QyEeokKyYI3scvTTZUMFDo4AhV8c2Oz6EUMKUcEr5j9WC64sOZX0x8Cu05fg9OFEXg0XaJE
Sql7jeiZb9PtnCeoCW6Z2P7VD4GbRDV1UgxzO1mfN1dJqxqDgT8Q0vWDQ4BF6dYEEfyT8iw3xFV3
4efQFBsLdUq81l5ZggqIVfq2MKS1oteaSPTmRrG7NfURCpVpoOqULTT0s3XJEXU/K+RBgyW01yMm
yLyvH1fjbSsI8460dIGxkpqG3M26QDBVtlhltshtN76T3tm6KhRcS4Ix9Z94R62pKeMe6NU5mi+j
4GgQDfve4O2V4HxmSyoFFDHX2jIMaKz+B93HGCJ078tQ+7uT0iXly6C0zyUT5cdRxlbP3i6hAEK3
A0B9O38EAchubKnTmIUESzpXjM1GTFr4eB7DUUiuRPOnbuPoc4OSVit/JgxmEWCZ2R4wR8KYx2J6
YNjfVxggm0+bASF0loCax5cbfi2iz7DZQsYlBngIp43Hob7U6QZB2Fnxt7V7qn+eJoeHjkI/npQX
FVrAXhvPdrJjUWIDYDgKOOHKdUchmamsEwpdbgg8PUgEAj5lnbj52Y+yBcz50+M+NdxMMElFvi42
lUPWmgZGtl/KhBcXoXJGLlWHdbBdbLKiaiHvabzYlHr/D8ez4aTU7htSPoof00sUN2RDorvoa6Hn
UWwnwq7JDIn6+uRnjvq4sSGO/PzeT6TNJ5tRDX4UYIC0iI0l8b146/ToPH0oXd2v1E/wcNBrJBUw
6JJD94BcyIQXh7pVk83lYCJj/JHdZHOWbb2cGh416CiXO3OM1c34I7HwoBDzhRvUuSRqfu69KN3t
wHccNTqgJ1aqAkapE847dVsIvmYqcyL2LKsvGu3khI/cVqzUFri9IJAL0kk5csxIn9wjqyvL04oE
gEFS1hgoV0OVaEtVanXgPtUumcFqoE15skaMnm6sNLv3A2OH91D8BNuG/gnuApkXJV/1uoIHFxTI
ueIRmQLaQ4IurJVqOFMT5Vz8H7e6q06TovwL27RbTQMTmS+bvzq44cOm1pGoY1vpP03sta0YDHKR
gng4fh3Yl9eZKQ1ZWMHFhC6fPL5CdxDidSVFhBgvSAD4SqrusKJVOnfLL38XlhpIzduy0yfT5Okg
gw4g314vVFf9a0hQ3EDEFjcEIlqVnw0vH/+TRPEOB6IAlOS4IdeCcO8s8+dc645oH+uZOw1iSPZp
OskTnNu/fpyOhKnW44R7WU1Zc7Y0k+dSWbgRcHDYDCg4dvBxl0ABoxZghjJ0q4TzerHV1T4M/94q
BR2iX57KCiswgtn3Nzyo65sILZbwa9maH8nUvG9ElXEayTfqCxrGmkYWrZSk0azQpa2GDLLApGxH
7VWfsPmUjpr9Y6hnX5RysszF223YQPJ9RSCfVSCf0T5miUEx65qJoe2pGZORpf0XB8obfLNHHF1P
X3gvE/PtD51fUI8uRiL7MoOfPM3BUvEUjupdNdyZXngiNmXtPL1LVZf2P8SH7q0vTo8jTj9sIAJ3
jmsZ7gp+amrWCnrPbjomrFTL/G99SAcCkaj6vs30ZtziFO/t30evNsb+qD1NbHcuD6invGTnfBnP
5SuAS5Kv6DdsnykeqlTacfacRoVa+dExXT2WS30yPkwv27C44RiUhUEJrF9Tfhrljc534P/AAUFR
+UYyaQ2dPGY9IO2xUyFTyf41qmLDOoFHSGbM/YnaXD0NNqbo4Vhj++Geq2YgiIW+d4zYnoVD8z9F
W85jx4x0lT5kB19/UDMHRVQ1MByTAgXLN7f0giN/TMA+b2G6a9eupYHMiyZ7e5bBFprgb2WduBxg
Kijlw5ubExLBjSCoFGDqgW0IjP8WqQHxAYK2yehlwbrQjSFcyNYo1CTcZEtr2eZomRZVCUw8eMU/
fI7x60eu+uEsM0C0GdozP4C/zdSpi/Q230XNq87WO2j3KLM4Fcj6d6RQZBui6sNmMZDfm6IVHOS5
ZxHdA9P4FBmVesYvTCYLYnWzcImYIcG3xnZfjWQ5IG9POnxffsOzVuO079kmMlt/bYYZHPKRzqAP
onO7tbovLgzHapEnitt1ae7q/e1ssiRZtlHgQdzUFUchp3uwEAz4KBoOXt+Ob+FLSF2s5z+spCMH
Qt/9md3Yj6DDyZWgDzj8wtffXA5y/QOW8RtBINIqBk+vjXkTVBZnh3TgzFvYq3FFOyd73DuRN4wS
ZDVOhVOb4Pdo1QN0QEO+mv9sOVFWIOvRsTqu4KiC9tiOaPpZX+aewa5/Z0CN4qrr2SU5K9KyxNEa
IWl9AL8N8NFVNzXFoRlbC4GYTEyi7ZS2t+iWAjnmMV9S0kzeiMGHjBDkGSrWa00nQNLrQuO/1har
vU7yGc7b2orTVyINdMGyyJf8lQncTQo31v4+vUCcEXb9hhUl0IBrnuj63o7qiVBwdXvBDSkDIexM
nk/GbWF16hli6Ke2qWKSA1k0eObqKsmLZ4m39PwqPcWiZv1SY5LkHrerc6IKUgsVWbW2uPbBR1sg
hkQejhO1pfCigWHHXtjtuUYMIDl2jXcpoPOlR1b8x1Vfqd87JejTuDWodDY3lrfXBpxKYlhaYy7/
6X38lIpk+o5LuXwkzJ+JbEZOKNf3uBsHJs1X7iHzP9/3Q4ZEyODC+7poSdMJ/oGO0mPvNiMMkoSK
lSBiM60KB+HULa+Nkm77JJQWYuO4YEHQedpzQxFNPZLjDNkKpVCLfurQJUX1BuAMkgBTYVebslUL
3C3xF1eNherQDPQLKazpZFWeF/rpz1SEM+PmsjGfcLcQpcf5h4y3oJQiMHpuFO1rnDQvVqcLogtn
PjOmyrKNbPVzRbJTD5lTb1E3ISom27DXuNxihiZIqlEvb6elHLM4QoPMEHf7JiqRrlj3PnnGuCEO
EuJllfoo+vX63CVkIEJhL10jFRb7udEk2+oQjrY7cFyYmoNQNSB6r6gLWRT6rTglpHwxG+wUfK+Y
bW7kSRq6omK/jKuO67h96tNrrcXG/a4ZqyJNFcdX6s3yyA5foYGuidBJbpB8UoCMX5DSM3L3CPk9
+Nkfw21601iqwlm1PGMA7BgQaBU9uZor+0R+7F55/Pwnr63TRBWJPqyyjMHT16DOcg7TebHMehQX
EDQKjC9hAMTb1xNWe3kQKx7s0d8QE0ZxuTPmDGKrQev3tn3raoQvR4/+8T0NdPOHwXu1wF6iXIVk
TLrQzlhA7eRUJvxWuGJ/q9Zxqm2i9sQr8Ys6yT8lEy+jOCtK86L3Wr5wE7qRRwqE1nWFTR0DNnQi
wP7Dqzi1zuWSLNpEmmjxMuPQFVqrZyLHDS4ptAf5nv8oTQ2Ts6wUjeW+cNjGtlqZOEGAjNS8tDt8
WlUE3vAiBNt071WgoZVrv4/6T0UDDAzpapPYu76CoM/FrBo9OvWrgXJJuPAv95RTLTeZ4bSGBUa6
QbSpYIm9G3EnZd9N2AaEDUwGm4Mw7P37EsqCFCFLzCsbUBNNIqKJJ/8Vr59LXUe2tjvTYY7SYE77
qPULxlKNS2pjg3CkLJAhFcFWa2FjNFDRqxIDzFdCMPCy/aabQQJ5Q+fltIMfJ8b7SgbfVfCONRac
hNFeTtL134Nn/PqIPhk6TcFx0BJUpXFSRJGnghLq+1iQrf+2GVZcxWn9J/tnYDX1Te+C8sIaWyKR
ioIPGMxndrypFLpvTUcGHn4CwRqjk757CpRcsJRp21xRxcRtjQZKpD40Ka0EXXorJiEQx+inZ+xj
fhTdZU55T09YlYqNupAJcvU/yijt9ZjzTrzg+7gEhTwab+SMUVxEPKk2aWMX0td04BOT5OKXfjAb
8me89IxHbEDVuW4qNVNzdOGT31OY8Rf9h5GbOn0F5At8904t5TncxeAoHLQrP29vqY6Km4EFjBCf
Azvvqpz4z94EcS3OUXpF/PiM3MJ0TBP8Q3Vfzrcik8HviW/rGuBZ1l0pkgPrvuJ/EIUNcmmpvlxO
3hzFqYsZO9h1Uub4pBCVqR8X9ZlOqSW5v0I43K3Yuy8pw/4Cw4QuwgNw4T0FoF1FCGmsfhFV9xyw
pEge70V2TEmpPPpNy77K0XP4B4u5me5frXchGUltNzxR2blZyg9bxTDxLg4a8qfhGPNHplAw5vaE
CjocYN3xhBg6e+vS1KcLf/YIVEJdWhVU/3BtCEBgezIAt4Nb+lbslmpKqVlD3k5J+bZJg3OSKYrx
ifSBVB98AwUoIzi2341uI9EcHpCImHBqCKfm8KmrK8qEC2++4R6jdk/ok2jQJP/qnln8kClccK12
eLaP6DfLcsx/SpYe9PSMlHQjMTYREs/UmDCR76J8ncC2ixVnow/tn4PESUv/LD3M4cd3btzisAfL
Wr60mg1UzWr7ZqAjQm6Q1PTNfV0HkRxw7Rk11Uc3n0UHmiPncbPNpu3mZkLipvYlxGhDxyTPfqYj
CQU8hEWn7I4OVlOmC6ovly4qjUbbUzZPL+SdoMf0rZs3aixeGU1sbhNpRx1VKSTeGSXxGKBui2Xl
6n2h61lGu7KAKjL6Jas7SGQMu1EXn4asiT7WNlewP1qzHgF/ek218CWcLEdTfKrhZ19wK5IHwORM
Kzssn7C5jIB9IMwzeD18gYOJYWuAt944n848pYOXz/hAfhcsNbNFvVkLX4DXaCBJbQ75sw5kxYlU
OUEO5LiSpOFBW/I5qLWmnRPtyBuAcw8xZhW2UBM5YNNXBQxuPrq4fpGhtri5yKyv7WUkhn1MqfQU
a8mFzbpyFVHFwN14Low24Y4KOmXA6hGg7cBV+Kg8CmlHTMu719cXXoINikmVaYVEkq5SC6HGuHhM
q748RsoP3UCtuka2GrtMpsrN0+HOww+HucWkiwHv5weuqYRZiTLtbSFCQZtkIO6BOzVFDJb/JsAK
S6gHxQ2Q1lDxmLvOpxKI8hasCdoLYxyofThTmmZjV+yMNK/yvgjBPrOCqqgX36R79M5OJZDVQPne
138h/PG2kH/G25lqU4EYEk215vW+W3au0eStASFZeBhmkiDrmWtfMDrWnE8wrXhC+ZrppPXYTGYF
oyUnOHIS2uAZwszwSpjiQs/aZro8rkji80oTLJZ3BnSWD+o33le6SnBKuyBsBfoIqYkGeVDBXXxH
LfR6xT8KagAxWp2/Ifex/qkxKU0N0rzEYbvlzvUJDoGMnFcN5is6uHbuSe/ia2lFJQ5p0hwmun5w
5vq+utQK/MUDQ3Nvu1EEcTi/x7M9K3kv4ibyaeOYl+WJG3C3i6gm1ZkMmCwckvaiieFA9IjFjn1Q
HpCD/OI1sVg3aWRnHW+ghMiK1WuF/52pmfB+SN2XJ5yQpthLpKJgOblBiU+V+PZcHt3GY5v9lVip
RZ4uekiDMXlHXPfQCF6ihS59j2T7AMIlVixl75m4sRmAIYC0uPi4Iawzqa+td7lQSFSVvITis1BD
vOWrpzIF3McqxLO2TGGpBFxjuaO4mL2FFZiGD4elOQMEcRtnDxYq6YG02rS1PWrLw0qLjLQEQCCG
lzt+TMiv0JEWf58KctkjMd2E3nOil+wjycCUMgH6GL8oIxYNEunmBpohmacdCLgPGk0W7Dzcr67I
1Id6V9Mq0xAa42HIe3p/9xwjmo/AsjZy8HvIO3QuABndhyYiTXJl/p67q5yG8nW4XF7MHUF2x2Q2
Hsro182s0DUK+pS1LDuZIObXYMpc9ikUMmST2/PYVvsmZQX2Y/lMMIUeObmacmadx5ss5pTH4oLc
cpeqlIlNviDzwRc4bsst6jRblnFYovF8mIQ7dAOhByEqf8FwfPiBePbCBudeUbDKdu457EGmLUpM
LZYvRLSTVrE/91r5PFrfJycdGvJ7UW69Qo9GFfv8Tl7unC5U7e5/uOwawGOA3GHDLDOyXotg7hUb
2S5U+9PFbMMAu218oZpuWXwv/5M7Ykvg1zaB5gXoXwD+NBQNbZk8PHl0Y7slVeNsLGRoZl88G4lE
SCnSOIZukFgZDvu8jnYkN7vJcWqnxYTaXfFLkbxjGEytsPLfxhrd1MIYBaw+1tNm/Ug+MTkoB3+5
tcwKog9+gxnuqpdeqijN5unA864sXJimybOinx9QIbtR4XrJ2V+GnkM5pcSsWdByb3ThamGYu4Gh
ayIil5W2H0qH68IDKg8C2eAJfzvPhEmHNdlWJwCWlZSSiogLHPQIdTwGpimHFD8ABiKbvYIVzfzd
x4o4C2UsbRqaBKjBiMgqyTlu8NlHbKcM54VZe6PscuN8cXm1Qd0mMyyBvmlN+E2jVBvKq1fxk4vN
yndVi4GnU1oGwFmlWjROtMVs+Zl1vnJ3o3p/oEjOJUHDxbK3jNarcDFZfaWY8IhzW1v8kg0rWuiY
UANIip1J/NjDMSx1Z69BYlfCZ1cSHosYEWAFVOS9NT804B7Dd7gdIloYkOZaI5GnlbGVZrSRjKE9
L2UXy0STt5eH53d2uYpXufOmsakasIvX5Ca6hZtB74qXXc3mO0+3o6kol07tyJRG2dvxr1M+TfoC
LcJ7WH94v0r8GN/GM2pTyvR9mLvmoVx2NS1qcX9V+WZ/nRh+ezSRdkXBDnJWcB3hCYNlW6//fUlH
2c6UE7FVnIyN4qDeqQtY1yB9pXrqOq7TqcSttvxwHErNtJoqbd5YY4ZbJXL2mKRAmdstlKn5bfg5
dt/yCxpthaV9XGPRSpcKc1KgkrOBLEcDPLS0XBeQqseJltYFZk2Z7AhxQsRcMA9J8gw4Iukr60Yn
YzS3Y2WEg6OtwYE6d/5Wu3ABKQeM6Z509YigdwfXOdqpXc56duLsp8CdK+7qN1pephdEUZZLjZ5j
RW+1Gegs+4KCoWuozRR5pGmPb+yAmoQMmqWlPsy7CGM7A6ooznw3hWFZwkvdKO7pbnPqz2+MtEi9
QAkzuoYgxTv8XUF+Cl+vqvX2HlXWv2UGJZ7LRpk2BqgJZ6B+9T8bMhfJLTj9MxTehG2OGbIu4bNT
Gl1ICTtf4utUq4s/y1Nz1OOSOSGnKLGdCt+H+eAIpUkH33TAd7dVBSErbk3ty5O96xY2SXKvkDQB
D+6hZZOTQdEhrFsBJQ4AUn+N4hSTIlE+xIAe7f4LK7g9uPixUUwVOsYGPJnr0FdUvn75QkveLn1q
5JNVDpHcHGMFbpXCa4lsIgGPan48mH7sCr4chIq7J21ga4OZbTulvhhQnfp6ZUMDFmjQsL4p1Bbo
IQ7HNCewOJe8a/wFc83QDDdcR2BrY6ldKO+80U65fyM6Kv9eoDdAR5LYFCJrIV1UW6xUvnL7iJyP
b5twnGILG0WBRluadCwpKEMxnVayUe28r3Xx/Pq1rWwBnbdOlla5hAPg8HCtBA0Flt4pqnoKpTTa
4HvYasT928UWwnrWLSJRVLavzwkZZ47o7oSEebh34mQXjULvm0GJqXDv4vOl0DyA5YD68R/4WUrD
Au7b4NmbMLRv652SszXW8loUvRRXN7Y2lnwPpfLlupZtLGA/HOXs+BW9/jAIJ67ZVrg18eZwMfia
L6vY/gu0BcHfZwHS+lUXxVuqCIyf8NfHO981SpBB8lgCURlU7neNmN0NHXFtEM5+Ycl07CVAHq7g
7tabUA5xRUVapPnHxxPWlzUJWaDT8WRg5JZnxeeM5LrJd3L+EotWYnTX7Kr2KnzQ2lcz4VAvpuD0
S/N4tSkK86PrU46LJvLAmPMoFDbqRn4JFPwtCca74Bcf2f3g4pxPiRVF4rUDjkhQOCpZD/E4pdaY
zDkpvqQ4vzbke0rFtDufa2vEodkdIe03NYk2HCACkjmGTUbG1L63O1YEQKU6mFjWKsFbgasx87ji
Qd3cLP5AbTtxp7pvvfffWOcskD+aFC/Z8C3TdFmQdebhKbCro+dBXNTFeHNoCrSNUqKMjP5GIkHy
rdgqitxSlflB9/lVMFhgDoYhoy9jzhYd+lo9AV6pwjAP3KrRgCN5Rw3dlEwpLGeX70RaaUoBr8mM
S/TVOzyIa1nvUFUQWOWsl7N5OuQvBguZcG1QH3eU0Amf0D8EBs3rJvg5BpJvQEVA4ooIsLcmRNO4
lf0guXdoUiyfbzGVQLTEalKm9niSDJ0y6+oMxu8UjesiQBe6dIZu4zA3ZP/IbCejx6LBDiubh7VI
igOzVXEJcK6QawO6GXYfu8z54LYP3a0lIELouFWPhRZIBeQhwpIW6/JKCZL7+gQFzzy0+09hQHVT
ke1XtqiFBCWMAY2y876A578TKTyJZB5p3Vxkzz4r/fra7fPTMhfe4k15gB+YCQxBeBjsDy8+yMWc
uCxPsUDLsRwyVPBMxuGSpwo3g/YBwLpvjD9crujqPSWEvp03+0Ind2i04qDOy/fTE86qqx2Hbc9e
UfLJ4ob+4RtfUZ144PzzPmBWLmdWxN3nfbNvtH2lMO2pn7sZXBqCPpRZ6CITQ6zOHqA/Kd5GOsFE
E57ENuGG6ogh22DcR6eDSJS8/0a/TeTgenSdTN3HD51TlWXvlmu5ARySzp9jj2jykwkL1njGLWLE
lq12VdVhwQWITNl0+h5KsaHyD1R08noNuQhrWhmg6t2kwoHcayZ4Cl2zxe5+HLwE4k0w4OpRVFSi
x+0J3Fb4wBjaNBoNSug0zfJ6AQdNzRqfFuvleQhhfPC4mjBZVLYtATmIc1wJHlguXy2mW9BoQRBZ
FD0iNMz32X2U8Z5+XJEFKyqi2FnlDY57xaR3rFYTi7AG1a5T9yIvtG/mfjH5aG14HfwcncbZsJe6
lkfmACwdWossXDxlBG1dw6dwyqfCjVhRgW26rrYZm8rYyC8gfC0QgQ8x+uno3NBXDZFR9ST7a7RM
izIG4e7YtMGKnabwQJ9/OtBz8OUatjG8jhAWrerHIb1y6tTX+DiaryOhqRzvspa+XmX5OM6Dgjhz
bq5o2UHQ3WWOogfzJGKYA0ynIEdZBCrRRr6C2r+aAgTRvEpo+wddlDlvyjy7x5+aDaTtYxt+GYAE
baZtTkaTSw8/nYg2Gaebawc9rjjyqa07Eyd/5trITK0oKw8R486ZqY6OU1sCa+k59EU2mwzYsCHU
HvH0fL5TFEDo2+2Frwxi+NHPTj4MDENjIuOvLV3H4oaK068oac2k3UwkGwnjs6CLVjrJdL4WM3mx
c6hZT6mLC0Zh1cdrZI86E7AJKYSyJ3kq3wUgDV7pr4LaK4irIqRRc/WlSLM+oM3HLVkf11LzElGA
KXHlSlJ3W+vuXkPIDv58Pk5mGmpfA8cogCo6qAIa99IT5hUCcHts9VzQ0e35aFVqh834wh8xe+pO
/9xp4sqFSeuOlBMJN046lI4/HsTPIzA8tUKJyi0qXHz1lzT8HoqF1Aoe65AjA7xYNGTEzHt82VVY
8lZEWxMFLfgPX2jq1V8I9xBtJqFNxsYF2cLXNc0jbZPq2nqEmPJTpGrxvdIWz/AOFBIAj6hfmyO3
2DT6bD5ezIr+FetCf7ecH3RfOVYHflEGrMBzSj8pQ2tAh6ake7pGr//x8hZniao0iVnLJ8ltf37u
lO0V6xZ5gi2w0/YYgin6ROxzaH3kLHK+JWvqyWMY68UMRmY1A1Gv7bse6aI/bJxNZYk8Oj1FmTvE
2GjqeIpPjEGkoJmvJEH+LQlJ7Mfx12v0D/OSXC0FPRyL0GcYGmx0T1dpZQYMou9dpZZl+0SP+rTa
LCgjyVCo4rNME7afy+nfx22s/om+H3xgeh8GlGlPmoVM7ovsgQ9bpfWJ6zYE3f/U0jdRwY1g5WNh
jbBaSVOsD9LNlnfcVCh8cn8bX2tlowp/IbxULSwvbDKZP2gN4uVjPBb/XZ6Rkj0UtlrgakAiDxkU
aYIfbJ8/TgpG054p856lg/dF/aSy3NLxACkqWEATcLF3kMGY7sga+4VSk3qIKuBmUDRD6oZx9ogX
uQysgonMy71n9M4FRChz31IOG70uRtL6UH2rGOOUcKejN0bw14QyZ38YzsffN2zMOnoQlYM8s1bA
5eTRYWCJNPlb7FnnCFIjCvfGCxwj9yEJxGSqQGZaN/xx0N0qv5g1MlaSNs9ymnQh677KcBP1VeTk
WHdzzJ+3mcCPI81LxahLnJ8wZ2ebO3cfqG0TyPIqBNMOyuqhoiBlvy6SerCV1WsJv8g6VFkXazRq
wlwgHv4dh3uVBiznPLuX58N6bL478Ano6z3M3Bjb8XlGII3PrjVw9chs62wTBFwL1tnNvOlDUNqp
ILSHVI39mOG0Da7BWKfWhQHl+IEXTubAbx18rs842xb1yeElFPnbv2I/CC/gCkXQ98VJghx/taXY
pmCO/dA5pWeG8J/4fpWmNYmrusxF/9fFphWwxtQbrQmMWo8UAF1gClzB8SCqwLagOTylhmLYthu+
xu+3cvDoUekQEKdTS+JywZ8jztVCjPsQGw6Wldh8Ph+zgOXxM3PMK1IPjuby5U5mz532GK3X007h
SFEc3VLGjKNmVdWxbaIrHzxsMINQSo6VxweOSKRpBdpy96xke8vQWHOqp9b2kXfntIMNz5MiLXF6
X2fc3SYBPgmzLliA1jai9cXd1FtbK6O4N/fWqrpzKQfthoct++MjCDYNg447VIzhVDb0xeDKHdKN
DWhdxX7TP+WBffWeIpNfqoDTF6bEW9KlQ73WoYZG8vIoUQaMLAkhZ8ePglWUDh4++V8m+Ll0ppT2
5R+4loCsm3X1pOY09nG7et0HUdPenIxsudJcQqaK+CsPcr9r8OxsX6Vf0VkULM0U9qBT0Soyehrg
ecZaCs6v+mYvbCqQ6hEU7jXB5Uv6A7f+1eE4EtwDXE7s9wFk57UwZGIWIyVgsJWKzUaXrJ7+rjLp
n6XaKK7HBLnU2piJM0TutBEOkdFMeW4keg59jrgwVVJ/sMsL4VBMXKj/2CiunwStoPCKF+Cbko/z
09iiO7Fk0ywoH6vWfmh3t9Rlpm04SOGyJ6W1G7t+p80TH1jpxFLeN8vdE/x+s5z9jB9ol6rBs4uM
v5AfNsXUdmWTxQM1saRuW22bREe6glErv4RicyF61UgT4JSYBEsMgTDAwed7LQ6o1dRI7fmsxpiF
ULl5hYtVQgj8Dtf+OymKQ+fQB1wsAEPnJaZJf9clD4L4UhbQ4j4K13EhUoiONhDW3qM7+HcdW+qL
6BslLUS6j2YnghTvN0mgLl+LAdusF0llXemjFr7gVhmdIMSvCiX5Bol8R0S5NTLZJ9kF1+eJk9sa
Ulbbh5j1UfSBvAKDhTdR/25ms02zmqyoqD+v871LCEm7g1wegwkvz2YbMAvMcwHoupL9hbH6GEOE
ecow5A5FwlnpLyLtvt9wYpiItyYvWBL5s4zhxOLSdF2kANGIvJfV8c8q5iHfSWLicJUKbitlVF5b
1VN9kQeATPLC+NOMTwLrMaoLfTNnYY7lz8EoePyBDgDonsBGcu9Os13TUSYhaOeX6yX9aBhbLylb
MNR22h6a+tgUx/2Kze1ZIpnyHEsQGxtc+Gl/s5sebH55q5nxAuiYniWzlOoY77GUa0NkKZg7nPYV
xagCnKXGH5FgBi7Rz0o+8fyIGW1ZGlOUdYxRt+VUGhkEXWSRfXqlQg+Ifhks37vc1Gr1taLMdruS
+Vedy4Uy1jo9O2W4X755qn+bUYi73Wpsvyx0wg+SDPx/ICRR+USKqE+OYel32OHTB/+Rg2nKygEQ
3b5P2zw8/XBHn8AWK8dUBwMc3DxoYhVAC/E0mktQ4oq8x/KqsbYYoEqWkEk4k0vYKBeBeYGqaMEX
ZYzG7f/S4kr4YKjRmQ/3COWUnbcM6OgXIW5uALBdVCRGuc1Wc/3kOa1F8IKBfN5qi05oGmzhMgWi
IuLRpXUYnJYSg3NpZviuYDiuKZaHI58cHZXVv/JRxQVAxqxwXUtH22fXadIRPU/6gmaFlzKqY0CC
lFOkbO/Ab7LpTUTN8+/JBxtAs+1ePPPPPnAcq7GtbFwvCrDg3WHFkPM6nwjqLkFgoxsoWrb8myfE
NLfrrjhLKQZG4Q4gH9Tr4DDxZ7UwoGnRd7Ydbmfi+iMnsq3Cn2YPGS+2BwMzxhiX/dthUDmYQeuT
BL5gjRlHK3EclO/wwJ6z7H9dt22/uYuhoLBw7x8Pbw04nj3MsEWI6+awAC8On7SrGcZzNCqg8zjI
QlJXE16iIJsBLCxfx2kYzC043TvU3C3AsZdsVwst4fC5pyD1zPGXDB78z+zk05D0eqAj3eEc4w5A
UjAEOtEr0znWjMg7xwOHsHo544SJE9cqeIITyqJW9gP1AzofcIQ5qpqRXgI9ETbQ1RGeR0B3TjpS
vP07VlsqOvc2YFHB4N8d5bC9wbvhfQd/S2/loUeUNS4Vqcj4z1gqWAOzOMUUI2T67Q7GvIRMWPul
dgjDK21np8VnryoqiVFRM6PlsWItdtwmYMo55xV6asIoosaa7O5IIYOzW1y7aZPEVz6aawxT9tmJ
i9nIpOk540zJst0N3r8Egul+6DdZkyomOiIgm4zDHLO70+DdWXDFo4w/oJ7dhhMN9xeLj0riHUxd
JfLTX77ExqirA9q1riJYfJ70cJGf8pEh0ZZe88emj7WJDcMzQW1ioGVu16KL6Q23eqU9QycXtCmr
pvx5/eoEP6cQ5dwFnNkQ5a+Iax0zfg6uM8U9wocMisEDHili9oudoHz5AF8RoW4VlDY/agxQtm8E
998r9ID/P//5k/UxO+XFy68PnRF2rB0jziyvvJGK4N3tnkRAiceLTRzi3KGH+BkL74FphrsFo4XB
mGXoCs2vC9Iex9FANWF3dQ2rBCRJnR1XqkLUFi4QXtA9Wig5wNBcPpeKOHOuqmYJY+wva/cEbcho
CsFiheZECsxfeu/t9aueq2ryAv2zLLrpOeO0Mwd7zWM11XvZY3LPiqC3jAPa/5odxWv3U1vVjZh5
/YiuzsAT3rjKiZ6HQJwnQSeQor9HfsyJBMoVkmno3y4OqeFovTALSCdzlOvm7MASJ+rQbAAXhkPX
JVELAAgTw5K/wzmxDxyM8J5lN4BojBjk4XegM6zKkPFGARkq1KD2+7JhI/pJ0jZo5M7xXWfrqlfU
y8B8+mtTMX9iH/Bx1wyUPnP3P0I0JBh4JRePQNnijjYdqs4KIk/NsdPLiILWCcd1msfYvtRwrKGs
bWBJgv/SbQ7QIIJ3qdTLVJzNSkimh4+0he6BftHXN9uVX+/nIrG6UHeL64Wo9BUOgSkoWmwCHR7o
SBzRfw0msAM0hekFLfIc+4rxPiVDRmxLW+fESG3Io4sixOO79i79bntdQWVnViqx3B4y0Ufvis+X
dI5QQmMjJKLblo300WmluOpSh08wsAVdi6LsoQRBRI6+6Jf/0nNg1JIegIzO7Q+0fCQx/iKK0Qtg
Up399cC5l7apm9QtXVq33IEgGenMDgGypoheIUyPTO/LwB28ehb0yie5FdIk6yJvgHxn/irpeQwj
3sanxz9YG79mstL9KS4kxj+95j/dsz106C9g2xZNpnLgkgSdgqymCk947GHKYcEyXoZ1I+2FLbVr
v3hnWUZsCcRdqNqFww/q4mnXZNfyQD389hIvi0nS6UVm7MLTjl6NcWv+S6qlx5hRv617zWntMKo6
cpQydn+LuE0moFzLFLXrx1Qnc0jtd7SjAwpB7bTcOI0m3bqHUHS+Kg5QFuMXoF9rEwLKQPjwLSxo
ypqhLKacZEMhdRkGBfkyXVesLglEAzLW+uluZ6x9NMKkxITFT7+3lF81EFKIqAjNUR2E9MOeY+yT
si5IvI/kvo2nBCd/Ar16YZaT4cY1PbNrL1g37xLYN9ctz+QgZ4mZJCBNKq19H8JoSxEZZi9/cN94
Iuj+oM0YOoQGeYLxrAJVuUSHtA8k+VmQvBxRJh4USMYtL9qwhXaxxjjvHIp8pL6rnmtQflS6TcT9
zjJOrE+6GqsZRqU88d87rwHNhltvG/nJNJvyVwBL0gk3RqazBu2FbnS2kDvt+abjIbb7er8qcECx
cPn2qJ2AFYixF7UX6+Uu7bWGnfS8Uez8lenSlcIsSe4oVt9lKRFYv62idm2j5WJdSEXNzGHS210N
nu48w6DOZdO9Iv8D2Vdm5s+QMl2EG+4E60sEadxq+UElmN1mhLPmsrykr/ErpfxhCz3SOEPij2cU
UIlFSiNfVyrcM+nPql26Qgkb7U9pupcx25NFAV2r4gAiAnxlPgQ4U94OappT/gjqypk9AsWaiCuA
WNN1aLliPs0GaLgMIyfYMTMwq+b9pvqHrOdasZCu2DYkZmPDbdkNPg8+qC1J3Q2C0MKV+gU5EC5G
jC+isGdoSEO/54y82i4ZZa6f7HwiNYTmnZHmC6R0HK7yFyklgoU5vMXwS6BqbNkVTSEZDc42bHQe
MCV3Ot63wt+bCXG0aXMGPZ5Q8YsXDVl5mqFWyuxwx2CYuGklrKnfqCQ0y1VTLXI+veZH4qBDNKvr
bYqiMj/z9oyQ9r3ghDDZHqeoAOP9BGdwUhNXDTpmVjcJXi3g8dYkcIOoG71Ahcg90PfkLO2VtaTB
/UI/GObu4QhBLJs2CQD8bW+6YDtocWwXELS/ww2ldd0k+8bYEff2p8MmhPxA30CL2r9+8ZhngUvQ
JoJ73XMFwtMdMq9PFTVWyqZvuEOzoE8ru9BxrvZCK0/+VJPIZMPbbwOJKlrHjWWKKcC9cVGFTL+O
/UaBXzBXX8U1vvfeP2Y9QVzZiZqFX8lAHbSRbnAd7kbuVQ6Zq71Ez58/CyaX0dy9olj0G0tckPjL
YFwFkjTuPC6V7XVzW8RLzmW1WyZev/Y3LtRq82T1lIa9OQjPKhQRuCtDQ9UE0O+cAPQgsDSDQZfT
FTR2Ji7Kiox4vh5MLUEyNv85bq2UyaC9F/RndCtEjPI+vPz7+2qfnqXCL9lWpg4UPq8lQ+8XJvKT
1F9cW5KqklJLOcYqxK5jbbJFbdFQhsRGr2M4ESNM+c8dOTCt5QmE/sdmGCh5/2JpW02ZWeGPr5JN
iJJ5vvpwla/eZ3XrIw4l0DVApYxu+E72e0ewzeTOkkR9K9Pu+DoCHPCIl0LradIr97FyfXGLJQv7
R4AGI660c0bNTa67yBUEWnM+eDFooyurkhtgRltzHRHJcSipz4GHgUKmVX6/LaQktwjMzv+0hTXe
VvleHbuDAb9EETsYbTxOoTasrRGJcvA4fqHReihidytPdF3MWihFWevVDNO8jaVQad82fICBL3Zb
6MtwLvbK8COT9r1QcQXDkMU1/2lIeHwGTS3VsxqxHU04CQOY7be/1UAmOttYZS6HFeviLVXvLkle
PXatXMiMDM9pTMdA6Go352K8g5RVVgBDdJLsG/c4UXLkLOVnbhvn83jBvPJ3POWoOhK5fxqIh9Ig
ls7sbE55Q2HsJRu8U0x1ExH+po8oTikqgbX63pJ912WnnKj2CgmpuBCR4+1HkDuuMYQbglgDt/Bf
elvXSHYd17VXQh8Mr0LW0M+T7y44tfjl5Ogwj0ywT2qNDeI4mESrhW8q39s6prgC+8F73JvvZJL4
I1tZll0boX7ZkT/teY+nAreWm9IUKNyPTWTWiY5jDLFoAtzv1wLciY6a870OYRPs1nmvS9MdQLr6
T1ZT7k/AYTvEk9ID0k5PuYhZIhMHDrPo2YVq1HWub+GmZQZf0AHY5XFFNh7jEERYJroSeUIrWnhw
sLgfZTzXNOg4MkrVO8ysFHGLXkJv+LEMXcwuR+ulSsmFyuYyv+BVlX2qxYCh/4mljiPrelQW8rhd
FCENjIzLWbGuOp2Orpv4asonewP/dMYbBzLgNJ5Va4GYqLTnZfvjkz+ygVfaywW5QufyWMDin6ed
G1T6bQEEFPw7aHTw2DD/J40a7lIigB8LjuyCJTqPxeAs29lgcrtivjlnGAIa3AArg/0Garqvo7D1
vCrjVLuPewbC6nyZteM56ipDo2nxlulegmOJA1YoHYfHg8AvEInKDvH763UiF6vEs8vRU0n5cfzn
pN6JHFHqgVtg0krIz8GbuIzzSjFSLYtYoQygLdzU4PWinRWEcjSh4DGyIbMZt4Z9SGQPg7e6ImuN
6e5zoDX+3YODeVIjnkrrskJkA6Gv3WVqqiwxqZ7V+tFNbmxyUbMX96AG/T9pW2gz8uKdYzraL1wI
06Z0oKueuEffjY1JgtLuKVvdbgWKIQyG53jJKNNWkBDVZoQTnH+XOcdfIKUAFzk+v4goKv8TtD56
nDiQDWqDo8e+zKBx2lExG7PhQbN2zUqBWKTIDhu/LFGo/Hk9MmU9uT3Lj3OLFa4RjciopjYIsUh1
glmIRYXHMMZGtbUqu2pEmWyYt+lbYdcr60+UaJmD4UZggPGheMlNrlqlj7vCMIQM7gy5ZnqHJPtM
D4JmGtLWloeb/Hr7Md/O3PFcLEsY1bQTR+1URAl5OluaWkmeljuQ+BL2125t7rvdyBXoMOEgQo56
uNAEAvtUp75gI6POwM2ClHjg29HcGj/7Fw0cpJi+hH9UifdBtZTZGR/RuNbgEf7oqhgostf3le8Q
G0Y9KOj9foPcd763jriMgZkQTS+js3OkVDACXgniruzJ+YOsjkPPWgjPaqJyygwuUrYo7yPYHmJa
EKTLTRqRvlv+YjnC8YZJWncLECTreuY0FGb8aTP+JQclr2Qiulbmre59c3VEbTdTGRJfIhRRJuw6
nFM8yRlDqIjAOVgo8qTGg5z5oPB0KBpcOrTFfbA29jWDlHySIT9rKoN/LKcq8PgUPTA5v3VPzMBf
YTYV4V30Vq8ON2TYbfJL1nOzTWNJPg4l0+TJ812TyizPkutuvoxiJpFbJjfh+nKJaQdgxCif0UWh
fQU4h+KxMUq8cUvLI4IM2VnCz5tq/pGOh7v0MT28FG+ApWpQ5VVKcJzxyBoF/0kEsYlA+pUSZh38
X8rQL0c3JupBLKWn0euadY25l2ZKu4Z7c6c2Iv7q4FOGqlGv9zR7ZtukxeVqL80of6vZzncMPXRo
sVy4ObAWRLJpsKDwPP+4yIPxUN32UATE6UGIP3DEoM3sAWeWMfFfTtWjhJZAciqEI3hdTeUAFC2r
Dui/y9l4d7eQLKTdGdtEsoI6YLNdtRhdtnSQ49n+ukXWyF1VejbuQinfpqZRp++SdamSpdsBhWgk
SLhwZVIiopQGfEhsYjUxXCzqfQybijMJTTLXkF2lgVWRV/OffA5ciylSv2NQV1wKavG8Vbw9b5SK
cxk2fz+m53kpPq+0uNVizPku4c6PPPkz4AGjchwG5xomgd1X9r3syXczMSTjxV2SrZVwqLX+LjW7
22LEb0gVNBNMyWSVquoCTK2rURX9/isoCk4FWPmSScULFHQVXdXWsrUhJlTrvYNLShv8XYyu2Buq
FIKrDgpUvYrF9uPLL2Sc+mEWYAySN3ULjTSUnoZAEzj03iLTGveEzZp7C7pOa0gTLi7Cr6StFQ4E
E8ldT83xVZml4Lx9ZRkHbjHXqO2m2bfAErb+/koS9Acv12mmKEMaL2yeQ3eTO5GWltvl5zRStmwU
nDIGgsDr+bx4+bKF4H490pjvThg1S6AqIUN6tGGDvqvcSi5jsabBCjfAs64d3nLxGT72aMqwhhZF
FCr/dj0tAV70HtP6bwB9ltF/XettQtVCpywcCtzME1uvygySqQrxrT+me9Nw4DuNEwNLL11KTJZH
wORafFFKhBDCR2BQZdiqwaZ28BEsrBgyCpbs81Hrcm9sHSNH48GchjAbjHlu61OrnmkhEV2c7Ovu
Ujg0fEkknB0DQpFKhDwJw1DDhbJptixfNVUM1xZTcN4lARlpmy/HBwgaPZi3YqifU+nDCX34LxuO
o/3BCtAYBb4lCqKt1RL1gh0L0RgPdpYbJyVN1mBHmvh4LbNlTzhRi8MyH1/M1SZJ0ZKdeCqkQ6lN
Ok8FZcxYm+3UBVXaMoVDawVySNr6pdtM6S3nBy36wtD3OF0hmcS3qWyWh1pmA3ZDuDQlsH9wjTDE
jPxHqyajps4O2c1nqMcyi0JPJZtH8VElspSl1XrcuFP4KqguBHt7ZJdtwDi/scqDzgJWTx+BRgkH
4slTdA/fcz9S3SDikrw6QppeSVbh0WqlZjv+2xyXqtiLMuPc/Xhd/RB1vfJLyzp/q6Cqq42gqoT3
7T4RvrK1m2GEzTjpHcvypjEat7+ZcP62reYCFCACZNVdCZ+trLsdtu33SrxyzBSkkSdnitm5mtGb
zsh0dV9Hb0vZ0A4loetl7HUHtbAMavWl6QSI53LCBBJaipb+UP99m8Ni0qfSJdmF78+AdMqGenVR
TmolFgbGbpB2kGtVrUQaydXHNQbPjxIQXI4FkoBrz2mk/c1ikf2pF0awFx0nNNV4MNObtUeVzoo1
VlWQUae0XdYHlV+4hSDYbYBj2Cs2y5Xkp0ljqTw//G7TdINwxk6nebj/CVSC294KM7TG9WuYv7Wv
kzGk+KDrmMFiD6IpLkjOms/3LJD4ZSLZ7rwAE3dYgzSh6C4n2cIykHK4lz7uUJtMZKgjjHC8YTs6
jReYbCl2LMJ87U5W6tdcRpEPM0kfp82c8PmG2CpHy8sWBro1PQengzjwocwRf/VEVEaZm+X7/F/V
fHESsjYgKfycf7lRM10v2Y3y2D+TJVV8kZhf0Q0TXJzczIAzrhzgADcorG+sZr3S0M+umhH/aNnE
fclAJ20m+LxwEvlgx5ATJ/g2ZVzkJEbCkTiAVV1GfxO6C8XgMUJrFEMdPU0tnJG60oj0tQK0daGi
gmwFFAx7uaw6mrhVJGB9eoU7hjJ0uvxT7bre5yoriCgseRl4ofWv1qA29QQ3LKglw24qyFeASmUA
b6CVzibwoiOxbIBR5NvUEBwny9N5xNN1ohmMyYtaekymppU7tl2GoMfYUjB7UexKauhNh8NLfM4F
0JzuVceq5XDgRq7MmD8XWF1hvW1oTBp07tz5GZCO+Y9kaTJHDZu5/wbXqKO1iBENW16sY6W8QAqD
gjERt7VndP6GlWRJrTVW/MrFs0nspJ1fHwnQKUIA9tit5jq9hpuRcGRGW5BqjKwHKdRHJr8hq426
uZKqDMVvKvkHg+wM5Ptk2VeBgcKx4l9Y2N5WWLpVjO1HGfCpuEe4pESUJFJQHZOqlY+sHdVKR0Ki
cVwo6XE4ZT8Ax/iglfUJE0JAI4b0nentjrCMKKhN3T1qAGdtkXJwVC7/s9fSfOZVA5+6zU68lYGq
CuYHU3bRR4xJagpdKTt6fhQPNTxqXieTlUI9Xp592DxbESVTBsNhM1BRx2fDzmyBbwCfOts2K8QK
bcFooyKRmRfD1nK5ADnewvm0s4RshsG0gD+DIsfVctRrpXMUqJFQoNBvUeBRjCg+qUSpnrbfhCvI
2jPGi0TinvIKbF8WWljWu98gRbPxX6RElFEiSSdQOXXA+0phRonNGafoGtWJNMt9vBZjFeQsYJ5q
SBL45wCe/Ech7UOy/B37GWuRsI7O6wDy3LbJqSM77VLFGtWHZ1sCc7c03jnUT+BC3cu/ODhFtU4a
aobVh+RnqaaMaokkI5/c/ESw/BkYcJCY5aS7IRHK0tUbDfs+iQWIS03zObM0SQg/oFRmXtoVZSmI
NyyQvMkm0fpC+YUSsZSZgHTIBSD3MZCB1eA6YuaUG1bMWZp78grycAM7g0NnXeE45zPt+D8XE6s6
9vTI86NR1ru9qZiDWZ6YdeTAQbraZMTdOYJ77f01VKb9iMtzw3tKbiAbIZo181PdNrbY56VTlDcQ
c4mnt0fcacBXLWsyLYNzM6ar/1suweMZfir/7YZndvK0KqrJNNhxJNn+zLFBCTnIfSbHfs77V5nZ
t14LaPVPibldr44vlfz/X1bRgIz1vp9cWMSNasXJlEYY8vEqpOkUuyxMeMVnPGXtMHFwZ7E6M+yh
hYhTyON9Sy/Xru72kzDM2lofuXbvmojTCphrKytiPUk9DqMB94awBW5ZSsHeHEIhp/oPXVgQWZOS
LYzCLzarLH+hVIzmA8Y0yAMMi8HZ10LxUPY9X4JOUhshxx8A8zOIIEfKBLcDmcRS5kf1GOT70yPN
YvPQozCyQXMeQTvs/x0qNYST7OZU+5IQtTZZ0cEEKvAZrGGWnRBxSd/pZyuy9TOCf/zdcGL92BFy
igLPUyGzEvvbz0vwFGCmisZSufC/BOgG+sce/7raQNClbmlLaWvOciDXu4jG2JzfTxy4lkzUbwbf
8InUy/qI9TyOiJabAId0cAKTGnnP6lGy1ps30QCvXfQD7okqI0bN+QUlsKTwpK4p5z4PILbMIf6R
Af3bIy42S+GepltfkH/NuySHSQxDJXBCAQ15ZEoeRH0c2D/sVEhbiFxuGunNnKF3SL5yMgSLR990
m3Wz65EtBzLib++sNnXHkweQAsBcYYD6hZAryGlf7CuAJl8/9XfvwzNDukPAfzhyN2vFA0v+u3kI
zE9J7WOE1fDLkqK2m0GTRhKVs1m3dAuLMgBLEiUvEAWNc8ei19Nr9WlE9uOD1Gg1hmgWOdUdG5A0
SjDsCPcoNN5/1VEojnPdb7Vbnhc3DuxVZWCZehIq0herRZ2B4H0TJoKZ5NuIKexfQ4amhi094UrM
MlhD/lLj0Quq5pFsTikRL29lddX7nWy3DVzbcqh6mF+xlnHGuO5AP1dxwjtIDRmInlNvgRX1X1uT
vdItTk8fj9MFgYYzUyCaJFti/O59WMaxh0PB+9gWyXW2TT9Xsa+vT40tn6ZPSivYLJ1DRA80eVbu
neiwa8gkS8+tY5M8TLYihtqCLoyDGTk7KUm4sa2Nidn5qXeZnT5fHXF+lTZneE+PDfj0g5IcLOF7
rpn68EIyk9YBE4z9kE0bE6BewdSKZaYZEJccH85HH50yZ8TKjflN802TZYyQdi9agrbwI1FUFcr3
QxqwGcUteI4xU1Iahfvozdlc3q0YJGtyo9BSIp3PiYrL4SIgfH2x5mpEflv0/9RwXLJE6YJbS7QM
t9AQUyp+F5/9mzEpAKtqTKSRx6Mi3KWu47gWkeZmkSSplG2NGSjriXnu7idlKZMGX1EWPmfC9Sur
U5nMoAm/NU2Sjt3p+wd1fWQLdoYyivyFWwyBWzZVX3JSn9msBsY7vfv4Co3fU5SLqRUqMQYo2ehF
FhEXzqeHpT7Hl5sMxauLeup3aFKECXnuZanAUC3IPDqIrQ3GSFyARnPnVJvK87gZbLo9riK6j1Pp
pOm9ymwzGTNpIlhmXag88hxJgQL+Akb5LSh7JkHuieaN7ncVN9zolhp4K3L/laCGV22SUUOZIYsM
u2Add/TX2acYlwLmIW17b7rsxOXJk9QcHWRusnF+FbRdvcDrZ8IZFG5rl5szLbd5u+5I/J/nA8vS
awCIEXAR4409Ctbfl3vqaTwpmNV7pZ5rgNjtA3QelhfGmnWvjmeA1QCmrfSkl1ce92Nf1NQ4IROE
+N72zf+dAji8Q1eWnIPjE2g+3FJ0RiHoD1lMHznNLceWLpEzS/JGSY0d8br/wIfa86OAMEQL2GSt
o0VHAEQhoY1rEGrbhzwbbd6Ovk0ubdz2M2xE9bC98tR34T3NBXoSjwji1hBNiSL20UZ+gaWIZJFX
TYnpIX6N/FybPgIdftGyTfZxL1BUlr2WVbfUFsVmUvJCpy3C5zprGJlRjL60JhmgccwGJPtJOWl/
zLF8IOlErjELq7Vyb+TdVEk2VrLbUo2stfDmpx+ux4cmA8GJnegxv6ZJSV19uCNcHdmysJoEqQAQ
2jfxiJ1idKEKs/obVSV4G1zGoNnnbTPUcIPyb8vPJQUSX6s8rG1cem8n6EpbGYwjHpi6/IsD7sab
s9up3fLRJOi3X2AXr9Cb0J0btTXfGpBz2B2Y5RyGgqQEmvIqHxV3GB/84qbNqLcGpzSCeHKzy6gC
7+TDIyTEGgNN50r+aejitxsBiecvFG+zb01LGgPK52q5bp2MtlvGzuFTp73uh4kmn/BhGmrsqDUG
IzzXjMGf6MpRxrY11+Udmuvaw5W/U8Wmkte6/bkT8bJrhTCvfEevlqvUQD+vAThRUAfXnzrJl6IA
HcaabXSJkPeL1rP90WUxgUwsojyhzybS3y7F3+pg3u2QCSLkerHcPS4Z0m8Eyomiblc3uVRD292J
ASkzQ1H+PENe9zCB5mMtYbgmyTnU7RpVfeLxfAF6+G/sgOXlQ4PlYfRPRR2HEY3ibSwETQeQvfFJ
/X8MK79thjg8yZH4WrNQTckt3ISuw+5CsC+yGjl8etofjEaSFA27QEgHIcn3oGxXGKOuj++/H1D3
6aTPYtqtVJvwaB5iRL4HXK6gjl3pbY3rTDRLxQo006vhbhNkG9nfFEn31s8WlNEGjcCb8owhZNIx
/w1wjRI0xHF4T37nXS2uNCSm+INatut4xLDFe0I60n+9tnWw3k3jLQXWB6hSFUSe/rVISyQtP0IE
Jr1k0rK5YkJuDSFFC1IJeqVGXQgWywS+SkOdv5EX88NDfKPE7QMVtXQb6WxaNwREw5v+xGJUjutf
hSMFWophu/IfWKJQhql3uL/D2cnZ2yRv2+4XO6h0zHrjFmtDeJd7w6Cj0NPwFhFPm7Y5RghLa4M1
Xz8hY+bh5y95eVCOUAfsJh3lnwvQm8njllhDGcgQtWHiUTMMuQFH65yDpUhQzF2vWFGdzvhUVDR2
2qIRqqx+pn3+S/GxjRnk46ompPCyv49XMfoOmiEo6lI50vnwPG5sPzqC/RidKhbXXm+Vi28KdHTJ
8IVdRuLuRDaHmX//umI4s3pkBv9fW4Zysu70sMlkzzRk5Lp+Ra2XrmX18ZARdCHsGY5bD4oLZ288
kGCda5kTT51iCfICA72w6KKCAAqrRvHlA2jAAPYNRHS5FrM3z7SaXXoxQb1Qs1QWDwIf74Unmuar
LUAksKfmmHnnh5EvXClvCw1AgiP/M3KM7TiNNCd04s3iTqC3So/lx046+inDXmdR67Id074XCowm
Iy4MikwR54QSXK4kCLvDPXgAW1Af45hfqJpJz0lf8/vVy/aD/Pg7IBYvO4WnZMYzniEBK3xk+PGs
oEisp2q1IikUJPA6G7b1PDT6ndEiNxp6oqUjpz8pTNhNovLDqKekGoWAfKBJdK3l5QNdhrYN3C04
cBS3eIMCkNZWVCYSiBJXMZkaclcp1Uo0u+GGpG4mt1eYD/sjSTpMEqw2FY3ZRkuq+mqQ/vT5Se52
No/oenWmXoikc40P6ZK17PVFEQi2kxM9SrLsozQ5JrgDbxlcO8KzdvN3JZ1o941AaZVY/KLzdnXc
JC+KeMTsLwsWIHyxoQKbtjsHprlVgoAvMQvAM8wZzR8x5zEmY9EO2cEYkJET48zlMz/Acv+qfeO8
yCMVKe6BrmgfLA0xee9eM0Uxppa9GZv6IY4TcS8y1S/U93V+YV0QscFhxHEJHowr1vpu0a/beiRn
OAqSp7Gw1FCUe0qMNw6AFypNUR5TPo8AVaI0GG0GDVMh2MHQEjVE2IMHrRuz1n8DLRbdo804p0sL
e3icaxxGrdjoR+19x1x5qrhfkQ16InXbrEkdTHspDWVcJdtnzNM2PmzzcChUe2eJzwIYibTBJ8qr
N8hElpQBLQLqX3kkapWgGim7IPuFPapSfMdcnpFpycCLZqxBPxIliR5/ZwrL2e68jvYqQldhgAg6
J1JRXXbrvqheFcSvNHbehvxYdVhGKff7yiaaM3FVMzYX2zoBLK6rwd8W6DYHZVbFtCUKtfTReFUs
8rvnTzVUulfqtFmw1Pw/qO89tLo+wc7P7F68Q3F8i/O0vhwdSDDs0ZIKpwTa3HHnaTgnzkayPQpE
2A+cPTRvHAsiGdCoqdhxA0LvT+6ijDn2/j5fY366yi//sedSz1CVGLTxYSi0pvDeH2Kqff4VcPzY
585FSeEjgvDLV1kozzZgQA8zlyYmfi6scSEKu5KzvaDkD+4aToy7CuQrXAMUnTcj8lxHYmJfpt3I
ewV7mRhAD2JLNc7HEAhlU2SREYghA62z6umR/KV6S0ueepdjGkJnuhGa9rS5I+tPD0o9XCkG9NR2
Niad/7oL5jmCKI07OG2wJDS6euRyevWwvOjL0GAjcYYkL92DLtA76YxCls2bYiwsBMU3NY9+EpUz
+Icubs2vDv7oBtzhPWw4rygMbnsS6xpdX8MStHQzbfEPY9aDs6ATNyEUfKJcUV2QBVmgSjzP/xvw
K9dUh9UK2nGOgCK4ywaN7oKPwiRN0GHCo5MSHJJ66x/Jg2NWXpWMR2ab2J5M9WAOSNUGRIOZT7oA
kncYptz8zA3gMLha/nrDsD9N+3OcD3sWzHCzjlpBDuuKgCE9CCUcMXw11nTB3YC8s4T+o0Bw7GAz
T7HRoVT9AU5ZTqWmKVjw98sK/ZAKJkwu1+CI9BpTAo+8sk+8TAGl5sVv8HRvN9q4LijKTZVnl/wR
oglPswNWbHyFqdR/0J+i0RekpJEJSqYYGyWruF8+6aUg0WbG76Q9MpuAevtoFVHPtDT6QxfCJf79
JGlorOsk6s6bRl7MJAHuzWdQ4N/vTXL8a9rmriFbnN5wdQ8rkmC0ILK49EsvOCXX53m0bpKeTjNc
Si+1IoHSVbCROTN75NQwNQMRSaOLso6pnK2HAOVxlvJUQhDYm+qjTkhhj2QoZSgB1Rv4bhmFMoOv
bi0vLAQiGM25t30G7aO+Pz2EgnJAsTAWql0fblJaOO/+t2LnJSGT8dAyGbLHuXn8Se6UUOEcBLxs
heaFyF7awe+0ViDP55j8n5DwcXhMJ22ey+qvUtTDLK7OInR7D8Lrrzmcr41xPkcS3oV49W5B8Z5p
6sO38E5pLVzcVW61apy5AGR9Lm42Ierh5ctMxFXj1e5gzJ3YHktwmaTsrOpsR0XGY+ozlIUYbYoj
74p1rL43G86f7VDeFoEz3UOcAVyZnGkLKsJgnvv1w8e1rWdHdvFQNzm5crL+82pUPmU5hz2Lt8b1
dtwKkIR3Pe2awyMGPGXktCablcdYKEt0qH+bz/lYtI1pQcm1jik8uEwh0QpgLcYl5j1wHPq4v2hG
qAXnN2ZueeXHr9eYBxrZvvJmPCD0ySwOkaPvEdPSoOLj6rbIcECLJAlwbUwpOEsGZAF8nTECqEaD
dDt/25tQLkqAz/wLQaSQd87mf2228R43QIIut+lUPgiK9GNh6MxSXn2VjQNUP06be9LI5erDuxhb
9wh9GelBh07Nj8wbZ9YwrD7XP8601fI9DgwEOI32jVNdJw9VV+ZxVYkOrxMMUYFP/JAT3GD+E4RV
zOU/++Dzlhs4CGN9m5ApgPmZFym2n51b5myq2CAPYmIKuBEkW2pa+ivh+gV+T3rVWiqg7hAJ3ZR8
6xWPkVvO6Ecjp+l6bUDfvmRlir3SwYEbd3y8HsnSVfgijXyWLlbd4G/tdXzow49Jh5Hen6fXSsk8
ftzaK3ZaRFtF0npbmeDkNSIEI0iSG74X7hVN/dYZpvGr0ZfffrLvcACd6chVQTGyuGd7byNCIHQh
ir97lQ8gZjPsLqUbHxMSZ/lUGi3Dd1j8nTYO83ZeJHQPtrC7wKRqKTxqaHVGACzDLhvvPMwzeHBL
Z2mPThOjJk7WHP11frzQZLnmN0wvjZbSVlPOV1U7NB83qvcw4jb+9fZJZjn0NBUFfrUFmezqHUio
76ajxCo+CphFvjpkDsobQWJcSAs/+uz/oSMYGyR2NyLpV5vdf9WD1HIOJNikiAiZkSsyrQgt0C9g
fBqrIGYwbtagPUn1tdOxn4ul3ICSXa13CmupONQCAIbc9AzpGDMKvhet2IgJgkH/FpZKJJCBJ/Xy
yeSvWEfJtyiWiKRle/y4ISC0dT2n7v8g6bVoNchIhWspYRvQ8PLS6+W5pSSeJF+8j2GpygklSx05
3MJ7VfPx2PVWDmduCPYd7V2G9H6bn8ZT6PnAw2zzOHySbJ31pYErVu9vgRIQ0JrVZJhqsI9KMzg/
J7ceALGUVtbVGkulmV9daXDGkC10GatQQy+NjdSFU7dI29eQzW47Db31kTyBZzrmWwdIdQ7kU/0p
vlEqL5EYlzWkbPpQ6bWYp88snjJzpDIQhEmsGahXiZfv9EWkuZqNmCqIaE/D4y/feiQPum50cXcX
BWM5v/wN+bWuNqe6wkMAGcDGGtkuNfVfIbRivmWrVBqlZy1Q5/vbEvmJQOPI5oH8JZAobO6LIaVJ
V6efkdXUnoPzbK5S1QipkittHy6MXeTTaGYgYqCLbsHTZ6M3KViB5MIn8I1U5uNgziZesZBHPGpB
LG4Yh/5g0UTHfm/1U5CGIV4uJlrfyjues8LtP4t1vOTk/MStYk9PDfkpuh9pFByZDTPD44VMawoi
tSyraesl6qo03ouuqY5jOY1pO3/Ifua9A9CviYK79GPOhP8XiXnIY9Thtt6NcafWJFgx2kP+hqrH
FZxo+B9D1O5TzHuIYBfGrxezsRoAIbktT5gw8aU1TQ3eIY8hixXCK6ZyJEPMJJMJQu2H5XYkYq4S
CQ2/yB+kULkgKH2+5imZBPk8UCtGcDlysKLuTpzWaCTJyIoeOkiJ177wOnbNx5yfeYidhUCFNLFL
1RT1bvf8vIHidqygtf2SPPa7TIE/KBFfgYxej6kv0uLuFsUPzHKoCPjvkTr1/vaj329uV196HjC7
5cBs6XAgiesDLjXeoaPVaiPzbiAyrXRaiF3OBFN7l/+AZbf5DDqoKM0X0QupxH2Bacw2vXazLs79
Z8i++FRCwtUKbd6YKqgvgWeiZHxBIzHWlY98mVls3+oUOy1OpyRSJlYfsJJ0gl3nTSNx5DmWVLSD
ga/jgEGHuhvxG8j0Z5zsqe0tjo4Zg3jVb+nRiwjOI6gKyFA1pa66AEpPLZGy/UO1wS/oq5p49gbU
71H44rk00i9AIPMUf6oom+Goj6YEYRoVye2A8p/d+CkBjS73gfGvaFbPZRfOVj5ndkkNVgQdxc6u
KawBz8Y/v3B6t7thr2k5PQzkaE4EjMW/adHQBZwt4verjCgXisDhuAhcKwTIpUnheJrxOSd364ze
q/JkeijZbxNPSSTiNAB0h7GIJY0IUlO9VuusPBusdawBaR1Yd1/i2VhyQtj0jpnulrwqoV8CEPgR
pZP72hHut/bEE2KzjDKjMf3GqzfshlquwHQAgsdZODJ6kDhWf/+er5S+KnwtI5vPAhmdnk0SHhdm
fLrkDK4ZCiBrnBXb0OJILQY02PRoQ5PTNumpGXnfcc4fBSBNchZPsvNGx+hpjWq2nRTeXPP3oajU
AzIbYRh7cBXBmR5H4foTCZu5CbIUTcqaKcj06hObWp/ApG5sg2GDGCbIDK8K10nNEk+VN3phoCB9
ft3vBNd2ckFfR/RJ1U9ZswrPxQO9KHQ9r+OOT4GDjPzZVKbrmHuSStFVNeFASFMSypwsdLpQweJQ
GOo5ayMQNmWoWvAjiXgAPrwuI1fRtkd5bp/amK3QoaXnXOzrxaznOPFbQqTFfSm0rA60AdCljsTr
OpgCw3bWAkKIiFnxEVAIfKZiRMyI5lsSCdYgoALSFvxos4I6bG1igu2MZbar69wZWyEDJVQ0KLdO
nQvAkwNc7Wc7mijpdxaUms1M3Cx0esjqu4UPf2QkoalrMD4LG8Sv699PTZrZLdKQ+8+5pBqXwny8
VBZOmi8tq2Tlf1C3eRkm48quhsVRE2Ubd68+WRWvx02r7Kh7ZLSHFPQmS6pWyonzRq5/+qTpJkHd
EqoafgeO2eghdil55Xst+tx9Tb+yhpZc+aMnOcfXe3H5/7/qdpuaJ9qxrKqqOE0vShHm96cGkXIp
eXI98plqZlCdlAB3gN9r4fNfyV6KZNlRN++FPlNh+PRuK7d5+lu2ssnGMfdsaOW66V25f8T8FPTE
SfHnVSVrphSuCdccKIBlnkjVdLsG0PLDnmismHmLvdhUat8tY2olMJrOSy/V1bufNJRG3sNDJU50
OIPVytZlkArNwhWym7I/Vr1Wn6ixOlsP4Orfyo/w7sT8i/uzI5092NTwSGZpolB7/DZK2/EQ7SKv
Ma/0wGYs2idCSPTGPnb0fnvHwK14GskI+JxYBvNvvKsgDA9DyVzxfO7oyziPsYiDvpri2mfpygku
2ngPNcO46BNlwID/ZlEyfP1Cxw8tXO9jVSagaJU11C75rWBKvu5KrMmmJSFiTVH9kHRMPfuDADv6
bHnItxoU4Wn6E1nG8cgOAeS14yMe3Tcw8GQ7uKm1fQTh/yEB8C8YVfucvJjwDYi6+hmXkcpz4FgX
6JAXp00rGicIc1Y2IW4dc42dQB0Wz32bv6JWwTyyLmRdEYfVeovogInvQAFjUahZqPk6C9syYwx9
0rTQsP9T2Onk2mMrtwRV62Dmr5tvaKKfb+h7deqA55SvY5WoHxleOnHPlSYhFdSRhlzRn1JjvkY+
f4AmrRjheMvmT3iPMVzb49nsLUWvMjLH9h9nndK+UVIbexwsLGgjsAp5XlYZPsnrNjR5EdrIwArQ
rw3KChKA5cJOGHZzGR2MCI041yDjUdYNOxYTLeevozWosrPp/MC3y/489Fgwjqc/kCEvzSG7hzPl
YmVNVqVx1D8cZtz5SPLtStHa2z72SNdybSYlIHKa8JSY4TtrgtKBffBOQWTZKYdz5/crvUfAWKd9
RqhpELINdob5zI6qSyoCvMPE0zVzH1JBdpCMZf6cJH9tN/AEaFWoohVHCpH0cPApkBmowd/oseiw
+MH6gnTwUak1sQzH1cQUOgaGMLVnyHL777Re+K94XF8sVnpy5JeNVEuiSaoZOsck38I2hx9gVZ0f
3Uz0pOTOX30V+ad3pShbWuGlpTp86f6cLOCQnPSkJYdB1DwGjD3SUdGgIX2yyC7FvMK73cReTsG7
8t9h4ePIYdEoTj0qpX7ztPUOAYCSzgmMm+GSaAn0k6fwVQJdBgkAs1PkAMDrJbcPB0uOYxAu0CTa
7hT0ssRxJL3TUWHJQbDnLDG5T1t8RHaL59+Ldblf+PLJ/GXbj0zz+wjnBP1r0lhhgm3wrqSBWCCR
qDNxQ747sXsuB/kWBrod/Kdh6mTf2sAc8k8IzSlJKrJUjZdtUsZhkZxxpaL29oJSLnrAtl/5fUa4
JUQA7B/IIDx3mMbeQVN5uB4CBcnI1hb1FkjNh76JwnEoDEygNsm/iT1ueOxhgJ2qmZbiJuuAWhGz
AOjJxSE8lPSglBsNzzZCgdWE+BQc+aKF6lfb53s9L6CBzDs8Xi4Oyt7O8olmmmhimTkF1W+JDOCE
gG77kuZSUuluu5XlF446qHdXVU3jtwDRxtejK+5wbrGnLlrEQ0k9YjH3yU1v2EBjbwnSWQHq3D2J
JjUSEnGVIEBVinIKLr4gOWo8UU4nf59T+kd5ob+5LFS2RsnQilKOS4DRZ+2YfJTgS4BvkuBDJvgf
aHCpU+Y32xJKmuIh0S9BlsOUCaqSIUQD1330npe5fijBpqm7EYkqQD9U464mOqVkQQeviYCe2m8Q
65CGvcsm/zqZvA+EJbqAb4/yBQgyLeeK1KAx75mkdlZCd+PECxb9WkbHi1p66/zNxeWKkV+9l35+
suU9YAdWYDpWv4Lsa/tHc3eKozeXC0zS5JOUvHGgExmA8/FjywvpWgqq8Z6Iw8yRJE6Tgo7aiqtW
lNmUixHyXy25V20FRl8KoTnaf3MW1ZAKqOZt9pLgogkIa3CmTSweHfHNTXW8RHTKRNZTnqeQx4aN
KYLD3zC+AeSvo1mjsh/qAMwaX+raBrlGXSaDwH0lfpEZavWJ7uQNONXea+kRq3dzDiuScugujAzq
PiPvzyX80v10V5DetpU/J6Kr23EnSqelj3wGl0biDhOyKysravAb0HfIgSHwVbcaygU/WK17ojnk
RZUqk8iCWJFOCXlNFUmRSMOW1KO1+OuuA5FCRdM36a9eLi3XZNdrB7uo/+MMdLTXeiQNyyeYgggG
Mxexq0394kkVSlC/IM9//eE5htoyONTTybeRzP6kD7A/3TIeJg8y3p8tSpEN5x/+fHaplN0IX540
PDYs+BYIXWSC99JVhAp3+PFa9pSdSU+LHFWunQGBe1huQxPOxcdVx+6tT3JxIP3Kl3EVK69bI5JE
0u75AOTjo80EKsvNogPz7keIlmFMM5fTrLEkQ0YYE5syahzhW3IKDKNajQhtQfViOOPJ3q2DuuPd
wz+ImZGQA1afMuNG9vumjAAogBlHGKwrzLpP9DiYYOx9AOWLg3t3UQQMD/zvQhvkhPqN68dX0yYg
sGux0KsN1uUKB+r3EBpHSipcsy+Jh8zJKmc1tGTeeClcmek8n2+4rrKWewA5QwsjHHBkOWqRZhoh
HZRy6/Mx013FMVfmTGXxadK8q3roIQ++m6cBjQjLdPOxACxzj8bQ2UteFv+ptHmfnwXu9Ju3MuE6
pMzoVJYEC2jjglAaa/s9rePVkHH0eR71gD/HodGjezEh88NxykJIgNNlK/WOAiZIdfe4gaekrtiu
QlOXm5J5oNLkEKbV1cZtZfP2LyN7UMKdvh8plEIDbpQQ6N8c7xaYeMpG2aYl89TC4r2Qt7VO1OmS
AgVoOsoOBotw9/CS020sWnyhGSe+rTzqcAxBtykSnHeOQWWuP9OvRqEp6wYYZXzBEjeWUyB27o1O
SYrv3Kxvovzfq055krypkXW3Jj693weMStiwz/L3ivG7ofvKoW2uf7A4fYjdyz9Omw+qyWGIdWj+
hcPHaZBLHzNXN782PpJxS9d8s+fCBfJYnyQR3+120lPQKvG7aFWQvREEwmHh3lndPzlj8UoK2m+a
rNActyFEtU8TVo+b57mo5wObnQ8vrXyYi3S1dC+PWFBRRs6wpYMmWvwejNsZaDlokzUDOsmd4DP4
uZoTx1U6M2xXYswMCCsCyI3fbHA4HA/9El8guxbl36ZsdbN1zEfkVWsb1JVBo9/oS8IBPrrTL9UU
tmppkMQ6joA0qKmWLtATZAO+FVCgRGTRKBAz4Sp/gexeR/ZzBeiYYYLcEb6GRV/Mpw5xsBv7QGU2
pXNqAvQb9alS7kTZe4VZoJnDqxggfcLGkmj8A5eeFnAKsBCXi1PrwhenBpCKlFPlmlo9mKDyyEEF
yUlUnpCpgw69mgBHJ//MGIU+jKmbkRj6L+618Zqso4pYB0Roj9E9Hve8EunG9QtfMniejO3Rr73e
FdonqHAl3Fs1h/ba3Vt6seQs66ZfBlgpN1WM1BsU/5QZ9O06ZZep6ajYPNQrZw54gzMOgGZxoFBk
xs7qtC4ul/4AwqLE+xDyp+WXu7wHWUT6v66AJGzdMdTVJjiXxQPR/woBmU/yr0cWWqCaXMQ0WeFq
RgbizuLQolvHE8Ff7OkEb7tPrbWpL35NpJwL9QOuI+SAQyF9Raie2N4HB7jqESQymepu353g3rGx
NFjJ8fgohcuxxzs8WpgNan+dmNXtMo+Tle7z/qbyJadc9NglLWeMutCTTEwjix0O/QGTgqI1fqP4
mX0sZc9RHS5tAphJ6EW23I3QkqF/pSGLtj5LCYdGHihs/rOQKdE+N9Pv5lpHmgHFW2DXLnyVKqYu
i8AZr2jbQLlamcxR1oDM4BHqlDLKj6s/RQrnFLkiVeL6GNj2PaBU9QQcAvmjio1XKzGduDtpHXSd
/Y1lVIRMGcHKGb6+iGVhgcd5cSBIC0oUvvyo8FiXnsrV6TqhzWPcaYw57lpndr77j80IQuKsYUnX
RS8Po23IpszrWRGQHxCZoRBTmYU/XJcPxlfks9MxRG5y9uBCVAb9tz8fU5BWam/rtHr/Fo6m8z4g
J8qrL1sCGY8/r8IzzaTSFGCGyLVBjHxv42lVss0FJF2uYKnzpnIfh6mphQ14H/yesfLIeifIZvD2
3iNq/oyJ1y7phU1R3pFMpTfUNgbPCfWMrpC9RtdN6ADRVelELNgQ/6ge4SCN9SoIRDt6A6+tpnhQ
ITC9VSc0Mu3RomU/xtdKdKLDa7L1fwEJpFNDyL0WERlYWnHE7R0aC6ssKCKQ7+qqgZTYjUBYIP+k
i21mj6jkr59l6W1M8RdfatYy/1Qc7DqHjUeBkI/AMesTGKbmFVs+I3E3WTXHULGs2LzbX5APImIL
7cBF3WE9xumfhUKCvhrd9Y8OxfMAUO33J9YtG4Dj63D5bT6hb8FWVha5XusQfvOlCbiBjJuMZxNK
kWuXfavGCKDcda/JpulZqCF+phblmFHi2jE+w1RSVVu4MBdx5sjR60M+8PQgoEQ9R5uj5JW1ZFPN
hyapcFETro/+gUvU1ari0uKZi+Jb9xRHEnhv9oVQnG6mq0BjnN6arebPyvEvGf8zWIcc+PZScfuI
Cl7BZ+stow5TG7VZIPaZIwd3GXFoeje4JyzjwS32QNGwd9kiN42pCCPtT8gB26L7spN61hMFiy9d
hDK0ttJ/ss1Of96R+1MSv142PoVDnhIKODJ07jC3unTz8vNzhC3826QzoABpaSdjhSA2uWUqC52N
vapwOZxmJHXhVAV+CQ6hFVZwrlc3y3YZVIfIh7ih+T9fLbmBa4jOVI4dw1HdQSXcT8JCc22ExpGf
7WEvLMECOXLEh5NmUGZ5OPR/by1PBzxAanFuza3Qdlwgac8yWDl/NeBO+uQt96Fei/w2cvzk2LhE
pfdBoceSLRaNwAETSZqUF+pzopl59PncPIJIOCtJcyFb38Xm7MhMDNN+/uKvmZGCiesNPf6XBiSi
NKFLfzYsc95fqD/7h+g3BVA74EGJhvNzeAB7pIo8IjXbkweUR56sxTAng0A0NfUGdd7kVMwvL1H9
CM/IvHAcPgyKCy1h/3MtzhtccI9vvE1/p/Sufh22OluRKwcfyEs61CdPj0eCYszsaT/oNXkXV8JO
ZO7ujk7FE3QWT2LQGZeJnANruUu7HkmkCOIbMWxceP1Pva0QavbqdnF+6b7Ro+xTwMYpztnc1Chr
fLazWcJwHy8VIbjW7AS12XQhQMSZFbtCQC2cRgv3rck5c3H4JwrD4kk4DRJmvYxw1WhUF5+JUhac
3r6xevCTTf4XmUA2n4dfZIb6UKAM2CwANSzwbwchXvWYCGizgKgDIH9csCNdoszosGbDGLaG9kQq
W+a3k2TQ0lYgrNb/pAKEhF5t1mBvdwadpywZtDvy+3o8GYkV1QTIp6yZhxhtimh5DOT1UQz4d66C
sOfUX4fUkdzPMnvdQklQlqr3iN5coYcKSWFlm46K0a1hlMFY8kTEeo0QtN5HyKS1ry6zHXmdhq+E
4c9WvVEgaoaNR+QuZUQmRKUs5WlJWgTZJjR1E0mweV/vDhFSrWNXv144CDhw7DHg5GHR4/oqq/4K
NG8t/6UwsMYSQGDaGktCRd8MaNcT2J+1/cZ0OqdOjIve92BYgA0YyzsO4pACGMoVAFfTqrWYEmSv
W0dpf2RDfdhOAExcisMROVekaEYocAX8q/lezHyHO/M1+ntBYYZWDIGl6ohQ5cMcuIEvOutXRqli
oo98gc7IossYUYFG+rj9+sfGqJ7eeWI52ldP7lJ8CJdu/BVo2sO7HDBIJA62ldOBMHuHJIg8Tos4
N+kSq+pplXGV2oeL+6Rt6W+QbSVJNfwKiDaJkzzdGME63zVgADIi0trXtJQ/K42YO0EQbyfxZGqL
0PTYJEPEOCzkpOXTADjn7Nz+xUHMHeN8nM4gTFCQnto8wPveMX3DgSPDhXNw7UTDuHh8qEOJy0Gk
rZnH0Uso/6uM7B8iwPTyPoZAq7EifZSPCiRJNXcOlO0MSU7ybEosUs5op/KHdjUS5IUSRmXU2oBf
4OtoutRFMowARm5PXDL4qmW6u7Z8RIN/Bq7tPIkvHVF8D/tU3jEr4MqGhUFkfn73r0XVE/lfL6+z
ZXXEWaQmbwUtDf39LZ8CdnrwJW0Rdm+CFra6CAeckkTrc0fI8Y5rTWIughnwX9wurbNNozVg6OcY
pkiLkuD9lBys2Tk1qfmOryhY3nrgC60amLMQbr12AT7JfKEkW996VQyZSNqlUArpIgnYTil6ozt1
qp5zJwiMqzW4/L2Zvmm7/bfvsIjKsABxh1ayyUgQSv5fhZVvZuUIbaMhsyO+t4g1WisZTPuIBQ84
dngBbVk26lM7SHOvKfJH30hK6zPwKXXjPLr9nVxKGKO3uGsXvLOyMo2TIP65bf+iv0oayVcp1CYN
ZH5MG8BOzqv3vmK1b/1ro5n2xDV5RAMtqD0uM4CCouf+3g5jpjStfLlUDFKuYtmeUV78RGzDU1jg
4ZgK1Zr3EKS/yeo8FCjxZJf3cMBrsGK5e8idfv6jMgBNY/BZMzjzGDZxBheTOKsWloBJJxKRmfWr
2gmJjqpbsnYhTq7tF6vMOv5c9zbauaZ+gU/SokdhVCZtnIqQn3gg36aqT0UjcVVZQSi72O7moPH2
bDAVfDV0VC7YcUKKJ+nc6ZhZcPU5MwbQkdP1PADKiyAi2Ln/aZhbe67c2KRelnFvDnYkdgSFs5sx
qOr3gUySG3rpznNzviUfgJZ8tz4XJwL4NdGjVXZ56zMiFyt+ScwsjGI5bE+uIJbFpbcHP6DmCGOp
b29Ive3prydAxVadkxdoSGMH4YBCVZJDfQagXvpE/mZ6xU8805kG89/TWEhHIxOmaIT+tw6Ce198
qrWIOv+L6nddbMx99SOIAZp59X4uE3F9TPcPwhtRH//Y9kq8qx2rAko/3MbXyeC0ExzjBwpOQXaG
67cykIdKxnPpqyIDSh6RUxkdNWjJfvspaUldR3ergZahGfmqzgBKl+BSsKce+nFYKsdcKWZ8UWG0
uEd7bsgyqpkdG5AofoOHG1gU1+8FtC3U/9b3DIM2wDff7+npbMODr4DGFU2DkvmcCaEQPrQQIOpt
22j+itOtJUWTGCqi7YQW6DtpLn4Vyhu4WvD8FziJ+IDeJpRevjvLldEA5JZyZuK5QwYFFJUU2+XX
HWnKdx5aCESR0ia1k0osM/Dtu3J5mAa6JP5U+rwzAT/uuSPJEa9B6QWVDXUn7YYUcgB8iImu1U4f
byYCW5Lc6p0EjxCVVwWIfMkGt06uOH5s0h7GR098JDODyGxdUexQugPefmDeFic/oMUW186RmChe
nKK2wnkiihMRgE7oUHw1gKlI9JMLo3+guk7iFwgBano7I+EndgBj70sC00hecFANww24U3gCrB5v
ExGNiFuJyGe7VggsUoLmRpFAfQ62SyDKphYZRJOXOznvON8HWTFhkiAD3vWiIcPtVETMhQ+uAPIG
xOyQwEcdEgjiXPJQrUeQM8uPQqVPdYI2Q5jrPrY5gUI4aB9o248XNNmlsA7aqMveLshIV8brqQHj
qY5StQkqRHLBVKOllzU6B4TFzd3k2P6DArkebjhUVj9NrMhHj4de1IyaWndPjDHYpb/lRckQ6W3w
e+Lv/D/hOTVQC/YYp1/Z9QKRinohVHCtza/vrb5uNlHqZVZ7pNMxPWYI8qM8vU9i97r4bHqwtdi4
rlI6SOexj0qEQIQ22z6QxgQqmIpWcvRizykeWpRniFI8hoLbJXPNwy8sfuld2ryV1/XEgsz7LMQW
nmGyfsCkcah+od3VNQthHgQagIh76yU4P4ROx8LICNRVPa6r3pdOXyna+FvqwDVW4fGNLT6gtj2F
bQgFUE1Pb3KYk4BsLW8AcwfaIBn3U0CyyC3cWUo+lofpAqOhzNjFXSU2D9J5eqlvv7AfCzOKgKe+
mNpLd2Hsb8G735FNvX0EdL3Qe6saIOfO6Y4AViHjLXxlH00mzSO+tK2Mr270IRzcBd3gppm9fB3L
5ywLZEsrbYWg+PW4cRx0pSxDtUEfRLeI4ljj3phM5OvGHAHHpQWR5lnfc1PqIDyC/bplPAuFE8BU
E9Eje2deqKI9pMtvmk7q1FLliplhvndcUKRFebEx4iCzbznRPmsToAx0QcmujIujuTs04AF3cqFz
HYB9Q++2RKaRgLDTYXAxEpgz3lyRzgp7162hFgfn4bmsO3r9golLyVqBtE8UiDXC1GeZ59JNxIpf
FVyGmWMH3evIqSKE1G0rxvO041iy1CUy8yfN1ojDSkSAYyoiubcwpWNxA3Wovmf97usaonSRFoBl
74a0hIxCwUz0cS3XALYOC5X+CYnZc9vCVYY1Wckdi7fKwbssCcXS9DVTSFIxFC/1FTOJ/OuT7nsD
FkuT8XcEkmLFBKX9BKouGbbH42ZCei7PZi/eM+ov7pJpasqb909QvKXj5uhiqcuI6US+BWzS2p/W
8Z4mdNfm3v5+vTMpxz6YF7YIgUluIjVStsZn13Pv9YjAyIl0wCG7vqij2CASBFSPru/AhqdDyFXU
uaunv3Bj6oT/8dWc+g3XMoJQawK7pcFkytKR/n+EywI8p336K8UdrQZe7aE7csuLcETRovEgz3Ez
z6VqEXbVymJSTtbMPQGeg7D8jiRADQV5ByglvSNEC3YvlrNyLhGOGVH8p7PL820HQxdKCJHdOSgR
KYiB5pqB2rvTuUFm+4j7ewos3yeXBjYLR/v/b0tVrsqGujx8/igU9i6zPfXLErBcbJdxwtvFHVPu
X84jAX5omSLwQkhAxlQL7dG7PLwhtE/0LXeWtPv9uKGsNICR892RTRsUukUs8AgfMHSgTTaNVe34
1a7ZqSvFjKrTszRoySXaRjYOwlE9fMi7/s3tzmwiN3MxNvFcT0DkaCGCT6HAARkrygdJc7lujxqm
goV3SCmb9U+rWFvlyRs4unXzyG8C1I/3CNVw2r8NO4pPzod6cyPZ1nadvDInTPPnr7Ez4Zr+LKlu
tQC2j80yZ/IR6gtCmt5anqkIvDa3N91bNRIbzj5Z3rWGYzxj1JKtNOogWGSehnGRi1q9wj99i0DJ
ubPl+fmPTBEBfrVgEktdIFW4BqBOIf7Vjw3RRfyiZKk+HMOCG00WZhFQrDcBo35MM2ux0cAY71DO
9TKbjSp4Q45uaBUB2YJ/wg8DSvfUD+ufnrJ/cPUM6TOHmljqACjTOS00ghFHxYBgEeugpqOEr/Sf
5si3dhC7YdeCWYAdR8zqYUD3byMUYNgN5TuytrGUuynoYq+yFchxQxnkiV0lLW10RM3trs4K+Ljx
LZ3tB6Eqma2Av/g9cD7GYesG0G2IUGuRHu+VkF14P57EZeGLWguOjZefe3gZPu4TmrhRYsAES3B7
b6Xt8PdXnps/LDKDsrk4Bfl4/kt+orUBRg96SIti4/6mOQonJ1zfXb3a3FZFUTxB72HSlUx85Thu
hdfFrHfYyqTwok5FkNxFcELb7HSK4o/obz0kV7Zywvzp/4+Oc7qRuuifiw7yr/H666NWuqhxZZRQ
bhiBaQ3SPZoYkkSTNSvo3zu5O5LFgckp9ISniZy4Bvb8Up6mqKDbYML6FKKrlmAc9E3NXCv185tb
XEG2ePkFLICvSoC6J3aejQ1C6i7ZTnRYWg6bT/3uLcywpGYYMaaYszusUeF09q0c120I+qgqwiKa
6werdfy6i2rYAFCCCUG2rCNaCRAMrRK9ALlN3qBplsRGHu96T5gRZjIf9sH63F+/h6hHy39LcsvR
+sBxGyd8Lc00IcBUriA5swRVPJQ6/d8ApBi+eLkXay9D7TziBPWF1BdK5Zo4VJlCIUxcrfSkvekf
ND+IA15leZp1JVNyY1uCPY7S1rX3uTI/gR+7zs1WpW5kCeLqcC4yKhHQDr7ruuRvoZ9zkwPJw/dP
8/WnBwt76CEd1ix6votyWyJs3/mc3WsqCnOPBlS84ogeWRikhrjGRBSk8XZFypAIZscS+mAVU2Qd
YEfJ+zhQjtnT/uJaSaElwgXrbrkaVzz8ZeVvmeEIzGB8V6gtb1s3IATd5rkW/xmWZMkRCMb8wvg/
jpxsHfPV/+/lUDYVulp68LtH3opEvBqetIDEEHrYxHkLoll8fwu9pXR1wn7bp5DTORK4wnrQ1u0e
REMKS95o5mGTdMhnpXF2I6KQBKg8bGcvwreFgxHHRXy+URjMspkwc8PvQwasjJ+Jg3jDZrvtkzcl
sC9kdDOmIBcEhvlPCzluseYkOwhtzfSZuyK3IHsypYxH99QEp4uH6Jlt8l6jX9SbDxIo835S6iKN
QN6hVnhgU2CagBIQOzDuKisTfhoEPPiFUmDIUeKiQ1MdXCePNv21ldM88D64wj+Q/mL6jLfHAAQh
DJ7tEb6XUbAPI2vjKJ2fECl3LjMJq4aFB1pX4i+PNDpoNhW+a+4cj/ZYxSxzL8FQd8vSqbMNQeNK
znqhjQQX50OEYVRF7+ByhKy5RUc1FbshRKEKSusa7RL8VkAmPVITLAspIi94FhlypyEkLolIuZP/
EuZI3ktBEUEfPpHo9fdFladpeiJsqkfYvdUJbZAi+KeDx+pawZ58znxu0KJGZq7d/NDAKtxYMKb8
G6IcN/Yf9PCCHUr06YZwEYoSLdkDol7D/X6a/woOiAAWhJ5vYMPmvhhMVgcFIxzZHBHyyl7qidrC
g2hodWVtTZMuaseJ7fDOz8EeRQPErvo0BmMwgOy+cKXdWDXcr/MfSnjOcvVwUjhz2y+CfEN9M9UM
A9FX43/buoQiwk84u/ij4wOrzrIKVIsk+3KQI+8Z18CNPEjXzPB2dxq+ckV6dKVXf7cIu4vXADu9
ql4xhcO8n7PkbMqGDBnFnND6WmyvA7CFZ/F9Cwaci3rQzaecDyfxzLiljflbw65J4MKtvB2RGUTM
3gj6NRq9gmIVzwPPflKfq/+zRpGZtEjGRVTf0JWrot3X3hVw93adPEVIO7Ft5fYV4+jbL5fjvS8K
FXeB0OtCaFbsiATuo5kKOlTkJm4rXvCcu8LXQN336dXlyCT9WAGzhDuSlbv2kOnT1Gr4RvfXEXlr
9dcmnlYIqU6moysmXmc3ir3wOHyaF0XlKV1qhL7Ijzn77SbP8z04GkaleTJ0Ux8F6ccvTnUXb6Jl
7/yhAE8a3UAFhzG/T5xORfgSXZMxqH4VEan6XUAb2/x4dVTnhEgGNC5op4jznPX1KiQQSkvqmjjd
FqY8k2eM3LVe0ZIQ35Hnd3/QfVuOAq7zAXeWNwhl7JGk1mSckT2WXrmzVS8MhvP+PjCQNTAGFzQs
jyohMn+QKtlpgQ/1dBFggJuJVituZlc2TSne9RIr+XZufRnhpbT730HtgpXc/+JyIVIboSdEAB2W
5V7jYPdQ7DgdKU/Oeyh/p3vblmhobq8aKzBX3n0Ij3h0PsMW/UBHlGjeLZ1sYOhEBccAfoO44jkh
F5tTcLAtdOf8hxsSkgVQMHXWiabYlSdC6yThv2gXjG/PfcneM2r8mkDDOk7IeZOGVM4VNakqmENC
1B1EgJy5Ts0JCA3R5sddWggtcEppojDZHgEGM3dsDlbCClNFbspWxQ5Lnu9kgqeAtphDs98Tee+x
7tMJI8KQYVqboVHetDR2mHWSgBxOoFX8DcEkQ0WvUUnKyHDth8TNMXsto79cY4vGAJ3fHsTcSfLT
Ef1VHgQNbAFXE6oR9Of8mXYoAo2tuwuV2eAesut/62WPM5u8BUizZjEG4CzgwL12/OSrPRkZhuzQ
NnNsTrD3qMHL+NJdjjW5jSwistHx3MQow9HUwnONzwqEchiGmwkAyDwQrooc09JYV+2m1dZUhd2t
1/5WBlaDOJ2eEeoel4fYOopzwbZAGL28JonmAB3p6K/sJ2ijLWaSb8e4ZqmOofP6gTST5TTpfZ6N
gA6zmJ7M1hY3EYPhOs2E5h9AVK/I7MyXNSglf3Xl0QT9AFmv+3f220topOU2CTXMCTGsALtROEO1
GHBfbVvEFd0o5vvB6TMb8XAYkCXFueVzVrk3EUZ5gpx/I8u2D1xOUEroZEuce9qDyU38hX6jMqdd
Gv97Phw9be93KNbPxh+k9d5YgWUku/t/UDcQOR4PRkxLpdg0EqejFt7+hpD9MMoKnlGgLT3qAaKS
Jv2Co4IgfwmcKJYfcZ37chq7jT5UbWLPUJjMZBiTBIOimE00Zt336NVetGTr4+TzgGcngjEbwxhz
ncLM2dV4DjLX3opxP/v1AmOqCBNWc1xDln2dPPr7Rjmer5P7inORrY83CsSVhslsudiN+oKgPWkh
jyFRXP8zrNkaz04M57+QbpRU69P+SImGQu421V4KGeunkRB8s6UVkzZafbaHSjxdD9R5VAT/k6m9
Z7up9H2odb+Go3L3P00UkPOVNWjJO6sIMiGp99F7xM/5QasoohPqme/5g1tR+5Atki/2rrmUIwp6
hf/3qokKiIhHZPohOZbQhRfxgNhOYENeL6KpV0v5nHrfmOtXGUT1326VaWpX3JMZW6Qfw9VQhTFb
6QzNoElghTxrmlbbXVGWLsd0kN61p0xaE4fmmb9yi7/uqPPBv68xtNvSD9sCXB8IOZ2N5wGeW3xk
E47VF2JJJVAlQUinpzPqQDaowru666UxY6Pg0r6NEkpsJl6RaVEiZ14pToVoLatchlrIwI73hZNq
/yirH33c30DYwIazHJsTx3GQYRNRfRsyiptlNT8hhVWOZRwvTlR1HmywSuySIcjJ7g1JWTVqH5Nq
aeL1N/l1KEU6O/LXpBz6NSsiNiDLCLmyW5qpNFwF2N+R3o1gJcCJPuHj6QsCbSGgc6AQ9p5z4E5U
w4zmNd/b/CE2pRSSNX/NkYFcSepS3vrzU9X/vWEn2QR2vZZUSvAB3zzW5Cxu0jwwRTSiB5/pgMyv
EVYOKSiu704c7O4lnyKf2J8EXOsSgALryb9UpM8rGR1e9NxksSqzmsiTjTNUWeftagz8V3iRAAuf
3eHY3Hfagen6PTKaL633IsPU8lW0FOBfePwHJtCf2j+HLWEFmOCF+kxbf5R9R0ynrH5T/QxjEQUi
uxF88D9mZsIm0ppzNsYcvX+un521AC09XCZ1Ozp2ehZjPTzBM7z8FjPKY4sEIjcRK0kxcPcqfVQ2
SKgYxSloMiWBdbj6cmO0z69n5EqlzsqNpv6agPrnXZOvwJl5YJIavliTW+q1BkqEHPwtkT/V61Ve
Zv027sECvN0dPmmCX0kplUQ3OUJ/Kl254gbaj/UX38yh8qtfG7iLfJb4mNKgyDZ83BDGLDo8/AvK
7WiFRmTT5bCTmnqCHjyRpi7ED8+M+PIx0SKIiEHqN12xSlDbhWYRbyPRu3bPTScpaLibHKM8F+pN
NcSv/W53fHOmL7RGRDMB8I2HloGsRHPKb7t6YOvwoTdYcY/qwDDwymyWsUaQ5D15C4eeVv000Ktk
E+Harg0AnYkxdWgrPL47eWgDmINcodt3u8aVxWwK7sNTV6Ggfz8I38mRKhEBj+yzgO35p5A1AP+e
T0vw7tgwsvyJg5944V4SuX43GwaLGOITetYVDkl7v1ocS9PHXm5pQBTmTYowte+4YEa8Wp1tg0uT
XfIYDjnBpL2YozjI3Jqbvfg22pqDENB2nvD4hm5XHkGIQqdVCerYL5MmVKgoEnKUD+/E/ynYzGK1
9pi9ZuEbuDk3psBTvFYCyahoR0d9RnR+aINv/ry/XWC4Qz4P73gy895iyhoKfL1+de24zZ7UlEuy
HFD9vozA3NDFf6mx8u7i2nm+WJZacRxMhH/BRBZafoVa2b0YyqlX71riNw2w4zfav+sqknG/VAnj
uhw5bafdIYZUc+Gmy8LAvGZ97bRwaFMCcVVqEW7VSY2Qiz5BklFUJoUZEHfWh5VX8I1iec6gS647
zsVV9kUOTq4T2IHTuIzItBWfCadzpP2zqqMPqGZ/xca7oaNvChh+W4SEzSn03wVCNp4WDiAws5HK
5zkea7u6UUDt5f8qV3d43iBdA6XGRV+oykOKzwdBfh9t5CP7LYNBIHOtwOemk/LlYcxC6zaEBsjr
yb2tH9nhyJcFn3+UcF1Fcc7q4usV9MmBv3TJnPhbaEzZWaPR9GCTfvBWQO+riCywRohkWuVk7gWJ
lWk2Yu64O2QTeeaZnp9qYkKeos01417csbmBmIYWt5DxVuR+yzoAessTMzJMeF1jKvceqxMUbZ4R
i2eopUQXoM50952Co21VAm7tJI/nPrL1VDHf40cmC1Y0QZKenH19WO5q7yu9s4nMDydU/WzFfxqX
Hhd6Oe9usajeLnhWy8E2NKpi34OTC1YbaZs8OMoWvmiSEOjkclKWNdwoDesuBLSwVlOBOWU23MnZ
t4yWjFhQyZ+niGqZq3BEs0VGyUz7dx4zPuwdg/2hGQ7AK3CQ9t4cTTTOxsJjyF92vDwmEFh6M04e
2ZNirorExcnzG93Rmr4HT0hJdp6+va2+4E1g9i5lLLFTtbbEa5AQXEoeSpjiC8TzDjTz1WzYufqv
VND1WrLsHhSpkOMh1vYnE6Vcv77/+BWQXxgOQtc+QBtFVSQ2H1q6xBhYgrmUc0iSK9H0F3BvHiBm
Ks2dajUuTYGGOKoduRO399WgebtnYGzI6vaRB7M2m7D8vbOYKdsuUtl2VHcX0runvgCcKoTOHEi2
VYmZ08JCvyzj5nai3eDNLZZhJyIp02erK2qho66BFkKljGDOMCnshKzt7OlNryvhoCTLxPbu2kas
WFM2owFb8OyftbL3xElhgFmhXbjkA+ELsTYORu0L15R67JcZyBjBMJds5enTMM4+l3o1baei9N+A
x6kQef/mgFP5W828bklMKX9C4j12oQBcJGtx5acNb1sD1R3XhEOHUJb+/LuVGqDHL8dEejlywee7
ZPT2LB/ep6Y5WmFzrV23CQQi698Gr7EaiOL+BCykZ0G1gLHS0//c0RIz68sBMti3XU0IUUXn4gKa
ApdVpioj+Gxi48Hrv0NN9w9NUncwmI5/RpVcFCXylJSOncI142qxF/P68SvSxjP7y3G98Zvo6zBd
NGWhGoaD9pnnBoZqjNPSeJyLNcy6echeaOCeoCGotJ1nKXRukP60GCOZmyeB9NnnebBL1KlQxO+J
LBE5+J2iTArgmZxpc1Re9jOlJ5TdgpAzWSLHRDAMw6xri+djhxcHVEahXiD8RkhdvmaR6cPMuQge
bjpsZgl8xEBxxPuW1GDRWWJxvfA2S+U7chiukwZZS+rmsO6fhkUiJm3Egdz5AyWPUuKHJtJwUvsw
3PdUyO+w+1k5+d7fq/Yc4avQw9kx3hcM06rzGCgCUl1tAHxBw/u7Oxx8Boe8VYvXDiwWSKGDjCgp
xFax1asrg5wO4X6cElaJiws4vl3OWZfDHFzfxrkhWhfSN3FnXobgK2TFvpNn12cE7VQ5wFOoD8Ni
+kyZjbbs4g0gKeeQOoYRe4fnF28sDBS2CTG0G+2CgH0Bo/AuHpy0Ee8AlyEqSxckSFBgsA7+21LS
1S8XKXPakv7LAkQ6Rw961FQOaVEUtKH73YWFf3f9kabVEowqt/KZAQ3PPFv7n2IBjALqgzxuxB7w
l9/+xMWLNPggF3KdrN3cST2ZsZA+9iJrqeQOIrLoMKjX3JpH2CjXrDJO4Hd6XXfZXnk3ndSJud4a
p0Tqql4Ygfv/DsHk6QHlOLtIVatV7D0ia2uW1tHf/LkU86TpfYfOjSiQgXfu2JQ0uFfthDphqO+T
UPPB0P5LpndYSCu94olbHP25+qJNhyp2M+wztObewRGQPBdqu7ZaT4hl+u77bAhXNY5H3zDckWY6
cLzhtJN+qQ2p3so80SkEOyH2trzqwlJgbrBmHcBLlEPZ74ImXB+dC9slxV3/J5NdImF4SjpPqksW
BTC1MBppY1cw1XrWUqfhIGbxw5xop7zkjiY3ZzmEsy0DZT6FkfzjjeI4CAxUxX5HzuWt/agbOaG8
hu4evIEOLopZESQt0dhYFVFGOCLfjdGS3VGD0RDWtKR5u7wJtrr81hAKIWgxUV07c8pwAAYK3pCS
wCW5wj+nAGqZzmYp2MCasHBkQjInqgy0I1vR9UCeL9J0LIJxswBEv86RZ7TA8pmLLQVfd2AswluG
FA1Z7tEpubiDPHt0awKS9IiNkKBNTOoNx7j/M3zsMzvrIOsceU7QeQVwY/emj+2kRxNyChwG0OoS
Q1t6cDxKo7UCzq9oed4oy60MxY5W9mFizPPlIPDhWb2/uZY3aBgEkJeZE+UWW605MxkE3BnbtVsw
a796doy+LGEQO71y61nJPyvRfOpkeNR9c6aTQ03xoKOFbVshGhrJZ0oUbrEJswVxg4soCzC4r7SO
39IJD1MoJmEjxQlL4P+gPMmLX8nGp6XgEI2Yad7FRLf9GLIFPS7yFzyra5swdD5g5tKge7rgAVB0
RgW6v+dSRF1kyv6rcjph/MOMcKxwgX6n0/9sBupmH/Dg/OLMC/y4MsiYaC6InLLDwgAUwqgGbLI4
OknlBVO30e8GVAKhYDGTCrqURMzqiv+MwgETOrwXc5/bF2yhxqn/csCOg3x/H+XcYLcYTLf0URKa
dQ9sI15F8MMubjS+KNx13VmbeyaK3zHNIMT26ab+084veuROABu4Y1V9tqF6m5p3JNJT3jm2G9x5
SG+c+HBVB+7P33cFYqv5qpl2ROuqTVqqjXo3wsRwV4l+JbKaye/VNAW5sYtb3MAghaoZlaZc/Lq7
A4aXvz8v1/cjHjY2vj0CmyGIDorvqxeYXqrkk4OUG3kRbeAvc/T3txgnQKEwsFlt9E/l+kQIb0dD
oI1oa+5oPvbCxjADVYAkB1WwHtElx802R11sO1NzwTCCG6Upqf9Hxwjh+sFs+Ls2BYDYQmAPb2hV
aIC94Ew4DWoNXooSMgWFCubyVUefZ8B5t3MDt6b9Fyck7btxnBFreFurwFgMNj/15sFf/gVtcRAM
lQpnM04jKYtvixGD/SpWH2EC9bv9xApYw4E1pKQ08ccVAY0Jje8gBHKPRq55C4ktSiiF9T5E+an2
83zpW/dFmF1ldShWrAEdctEfhGOoOeBXyXH9uUDktUUJlBMPfZUpYa+A2rKxS2Zs4qHVYL78aK81
pjwwBohacgHodPObeMvCStG8TuOQYHgT+pFyOydKYgaILpRWU8u250PUWKzsZ7164dkDh5Rt+Bej
CSoOtYncYAln2lShpC8rU3atFIir/jRGTi3lqu55XHnwtxWibOCIr53cgomNdOopvxPe7SwtmdsC
SoHvfYx447z4ptQTCyQTuRrp1/kRdGoCf5KjfznafkUwGJ6LSOnSvn0h63bTYvxoQIL4FwwAr3rr
7fi7ThkZmYYUKH0DUNpxbjjXZvqA9VfRmAfyuhZkY6uZdaqas4w0EbTzAi/K6wVQzx8OdKYaKV+V
fl0MEc/3mf7V+UtjmU4W34K5N/JmXqTGOKr9M+1euPnZmAzbly5oqsnm50LA93CCMXxfZDJ8BX/y
Ges8gGyKSJaIT85KzipmOJoyp/PVP3+jZ7/cCbId0biNj5c77Ew0LhvNTz0p883dzKjww4xLNlFj
ESEpxbqncLZvzD2nKdjUxKfDjFdUJYJCSoOQGHqvhDk0BwMOOyb6XgWw+KWjL08ODjEH+3f+nvLx
cvf4czwxShPWuFxdS+TzwbHcEPZcILX/QlZFzZ4PFHZPlrXJ632adJGyDL5nvNzvobggc22ML5gP
zDUhip5RQsSWCMPU3eHHdNe0ulAKMj5tXsXOqGd2+vcAH5olT+eRKcxJ5pcewhLDiynbiRoKVn5Y
hrJPT9pVIEZQMSTJd53rGVxZJC1N89ThSlkIEhwTxAdOvQZlpSGCegxmK/DAhv+VNqn4XbbRURr0
20LP9/BqF5/L5fV495ODhSIq0QszVv3CC7HSbjowoFn1/WVpSnhlxyuBq8hiuIpfEFfyQNllHCDM
K2FWIIH3sPS6IRDagr+EOkF1K/lxSr0IvMNNhid8QxJE+mCYY/NwJV3oUuC+CUqr2JsfTdeY1hsU
Wa5Fxzv877LBT4l+8sqfzFlUYgLY0YtgGh3K1CCRtVXzUjO5LfgvjltZmE1F0ECWc2Eom59iMh7t
9OOmHHMiUgY/+BkPdcg545IRTTfN7Y2r8JbUk0znkl3y3DQcA71ZlxyOLCTgRt06sD3wQhkz2tiN
YOAM/rraTYDsuML3Vd/lstFLFhWDLFnJf20gQhgaQZhkXmhEurP06suvXZUwX35tvFIv0uWBwXGi
s9f31o/USfE6Hl1smTJWE7dDW/uP+penIaoWrRWclhn4HRtmYijA/+haRD7h/LiqESlMP73pz5w3
JhTOSsNANGMHuBPLLos+TmBOVrV/72ElKf0eC7RGXUiS7oe09LcR3XxYk30FgvtM5Tu7+04x2pLI
RdUu8RbvQDSnd8tFQf/+mfWViPTJFBMhyk58OigLxBbeT4a/l3XLER2hsNRr+m6yxb8WyOhVWSqA
4nl8+wqn041ZgQiZQgI8YSI+i7uRYGb35095yI8G34c1VOTHP//xAX0WIp6wYb6GVh2AXkCYGSFA
GF5EvCVSSf2B070ss+bddK3IW98FKrX+0G2WAVq1xbKUMOjwEjEhdkt4KC2VpTxvI4HS3ueLIDnA
18rxJSUigjUKPGKMsLnkfjOaL/ZjOUbxsF20vu2JKK7JqPvQamErkNYx20v43laXeA/oIpkRzMpR
2NvTDAEKZ31mUpahIhaUrLm3vMX4FJpZ901I520V8iDsPGbNTSMa2HlC4vSgSe1FFMhGtWFcgz1x
3NN5ddZqme6LWM5Tp6zIT3z4Pyaho4shNLtOIlLztZ2yJflBvUIWJ8eZ/uED1f4TgKZDyszuELBr
+8ZSWwBmCxLIXa6lKn3v/s1VgodaJJc8EdLflDUymj4nXD1xUkYe68c4+JgaNSfJgZFsDi+lVQs3
qwBo8GkV/Hw3rKw4I2nrTmHavNlYXZXk15Tc0H/iBQtvGIkPGWPkVgUiHpVIsGZThhxb7+/6C3z1
+XJZL0taJ1q35x5jX2/nBK4a6LJ7fvd2YEES8CVBK16Dfh1cEJkXzJZVCZ+bIBZaUcxqEBn+8InA
koJ899XDHvsOsYOSeLYHLutUb+BSiy/2WapiQwedGhIRRNQCJfVYPr5+d2sYL2Gq77iN2blGIfeh
yl6Dx+BM/jgzBLPtkwN4SeCcnNWXCS9OCmWVYayDY/kKC0+Ndo8PzQ3cZYQpBMLk1ZukkdtczfgA
PkIaSsQyG3ZfQTUK5+wocvH31twNzL+idKDn8Ksr18amxqYqXm1FN3CATTMKGt8vbJTQfgjiIXSk
hb+sC8TBfxOt+dSUyvGMLZSZJiQsaAmP2BT0crPLvB1ijLpdSZcMQKZMEq52zSg3xlj1Vp8MwIY8
fAmDLM1UJ6892oHIwHcedjVWzcwctuFhL9Ha+f/V8aB8Hndf94zUDzdGbtS/tM4cutiMuZe4fonY
v9I64TKIrCZybMoApprzYaZ0omc66HAEyJY/Zz+5bmCI+fVimrAHr9TbVx9DG5ehWqPo84LxovmP
32NEZL3f9qeb3vHmlYcELgDWCHwK/VkhyAJ7KCB+QpHG7QmPq8wNtD8bqvwFy4veeX840V5UGMkk
nqHs/TXv6SvVo0IhFLAGiKi9/a8NuJurxjmlKA/GSbQFmCnyFuRAj6ErBcBZx4kQ5V+nhngfcXsy
gRj3qdKRK2Fu063+52TezC6qb9Com2rdfIlDeSnBYWPQPozIh6o1/ab6WDVFS58cokV25FeafOcz
a3HH+mVsPuH1paUfWeMhjbrCCesOKiT3k3+JU1bCudkUL3MOAxPEZ6J6x+405x7xHi0eNWJvrD5H
h1d9OBy6GbV9U9cPy69mxlyASKRNkDqVRCu5I0T2T9CGuJeB0K+w55aPrSvkpaib6squ6vhCj/vT
N4J/5iHerx20AY63Eslo6xwZJZrsDgbzZP9PgWZjFEjYSs5SxkZ1OUhq+RLvpb07/pBXuTOkoXzv
+bphYRX90mVR4vpyeKJoY8uaxfPpjGIWYpikbBGG8oF3j961xtNlg+P+6Y4ANyw/tQrBH++ATwg+
fz/+UEdk9UMoHl0l1Q7/sW8/Qsj5AfP/7CUCTHbQKeC9l3glYi6izEbQpNZHOOS3jAyB2quIHvn/
mo2p7zk950pS+fVSTn83LzxtjxOL7eXkhLEmIP9UwWGbgKcokwxS2o2TZcgn/iC2k/tEKMrcR03s
DEKTbJZRQU3Yy8Mm/Otmd4mEv5hjD7IVuNYDvb5zLfSfKEiVgp9KMIXe/jUy4H8jjys0GD2hCrnV
agtGyFPLrLPMbGYP+682S2jjqljJpFhXOobWbytiw9KL448urv1OTSyd09fQlUyJwYsGf48nK35w
qNF94yXvW+6q73E4Duuj//MEgPHPTUI7i/3UZTkaATnGE9OWhL3icfJSXo0CwK+JOBaPaFAzWGII
1nCnoo3FlqgKrFk4SZG+BbUh+BL4SxsGD2nJOLrCgx7AjnGEQvZah5CWZ3nNhYan5hQ+XteklN+6
Lat7TG1bc2R/yIYm6YlrRD9UPSbBn9xI7AfDOsbtv97BfyxeunHBii2kP9dqCGaw9r5dLCYGkn1I
zLGjyKPwBULlEARZVu9BWiqsJxn1Z5dsjRD5jNbnk3pYXxTyahpgR+5CeZKr58yxtSfmAJWAOfPN
IjADQKC+QWWpScv3Pi4bXX0QXWtPy5NYBrU29vQpjWUYdOA4Z43mtvhGdFeeci3ZUDGZBsfnThVZ
3M0ble0uQzG9RCLKx0RcmRUaZwvNqLUsciT7AwhUX5AHYz9NcHqyX4t0j5NHcm02GxdipdVq7S+i
J/tCOBasuCHAMrm5wb3xA7vGCaffx4e4zm9c9A4agdsjv0yz9NsYJ6ju5tCMLjr0t9+B37N3c66o
b+jKokIPZ2os/IH3i9yJLARirLeVpWYAL/Aom8rxgxl729hNFHyvOCSBxc+kQwbGi6zFAHKMJPeD
dcHopOQfF/g0BfpmHnHgY/eL6AkNblesvMh3zCQPixtxgsqhqOvVbGng3HXbM9D0ZhKWogwnPFb0
xs98H7irMtLne5x9hOmh6oucyYKtM3EwoSEmphRl7fOOhJcvRUeeLDdiOGKKcW0uU+YYsj/UEj75
H08XrX15xfECO2lVHXaiIk1Wj9rV8k7gGlG9SVtR4ptiUiRdJZMevrUJAJPvmRDk1I+bNdWiJ0kx
zs4OH26CkP0kgcB3Ic7ZmmiEaA+0DrazDM7dNO0crx/RrTPJueRcZEB8PFLs20umwnqwC0AIeuCB
4HiERNGs15/BV7m9frDdhW8ma/zOvGdekXP4ibiBEmr6Lo0TOBVDU2QEX1AzgUH4raUa5zL+k09a
8BVwjguPGQ7WcMO1PqflN9KnTEkXoT/HWe32ypdFjiqzjm8APiKtlddDKkIrcVQrMj4OiZTSV91S
6PhvRKDdbNIzezgxu+Q0lmd4tChXHakxTDoem2cLQHKzoHYsPwfXGzm1tNpHfgt10FszFvAVtb4U
DnoPTm9DprLbKJOArfuys9hx1JWAMJWxYDZzg9M19XvzTqFYy0+ibmADbNbIhIZvTEjMw58P9dBC
YAbgrcLCQZpR24i9V4Ypi8f53nqZ+EPkizaT6TkNof8zPxRia/YYk0oulvT/oNLm8xSC4EmDxE9q
7FvVqUJNVJnP93+mBqMT6Jl/R4qddGTECQ5oOWCiPUtm/V8QlAuICTV5tSxyIV21zPbl92bhk5ot
IEgonNdrmgBPR676WUseFx/oanZ6jQfareTTe9FEO0zbIvDNLXUl9yOOKIshbGknpZKHmgOR0VyM
VjjZpzGBfNR4C/YoHzRGb0PA03/xUtZ3Tqvk7JeETqnpUD7tDt6YP/6y48O5I3eIKyG2wUx5yloM
pE1X9pfx8mZs/tbMU/npyILgKqOnuTc/MObyMvnx9zn+9HV2RETlrF5aGwReNKsN17W7jp/qH9fW
lINdEzBaXO3MsRjAW1+smU16zWUp9DEftE7Xia7dMkAa4btFYnU3ZDJ/qPOqv+sR7eljLrcTnOSU
ugMC7hh0mFNJxDadAzanTqJdbVdbssc/fe78HdaVffK3CQhb2rnkDeapBQlW8OmQ95HBHbXUsW59
/49nmjKAqLN2KOaEj3QqZEHk3N7RlhFrwVqni4xgdqDAMAm5q4lmm+F5BAmjxcX6zKa4un64Ikhm
SJU2tbvjEmGOGvnneb5rirft8GjColmEp3HpYFnq6TQ2Lxqqykgfr2rfRpOjPdyniksDVNFzz3VU
JCJGoRqWCUln0NMHMW5dft1Ayz/VjBIzVshSJhmEYUjxvFTnE3pa1XUsPHYVXWZaoQybU/3kY2dr
hmsRSWTswPsDUrGzniyVH1Jksyv+RA70hLn2P2qnVmuqUmq8o/frVS0i3M9+pt0dRIUSkx4P7bFM
wXclq/MZoA585kA1k7/99Npkcb5jV8xXQOW0MJ07Sl7EX0BWO2QiEIttsjKs17xdj8aaCik6edHQ
lynsuAnImB8nRql/a8bbmMfsjYDvLE1Cvw1ddVgfi0474EsfKiNXsGWMaRjF5sx/jTQi//t+xEU5
ouEsP/OdXp8KpEfai7iQzJOa28sIsJNidoeJyG79bFfybUz4ZyXwxqej+a3zBf+ENLrsQm/DDZl0
V+Jbdb8AfUcvla12l2n/pfgh+sz66SDAoMbMbwEH7JOmv+bwkUPPGVRIq6M49sswkggoOwyBUNzA
2lz0fA426mr4dv1mcsTBzNo8q9Wm9SK5ellvVNzoWNuolOl8TKwzlJ/v4fg7a45BGSbITcWC15Qu
D3qyMX0IXXvgpxyPqnJCMVV+mMOrrFOI/KuBy/xp122/J/A/bBLU2nnxEg88QpdwGq4gB9vScjcg
UAMJP1vpPDg8Egvz+rsrdf+0LtUJSnHsey6QajI2lBaPJAoW63XhsuYrfNgnhfaMObcC7kAEQGDs
VE8FQdf9KWir77YiZkgxt03G5Of2NDBSjPkKXVA9BmAhSxG39T6dVXDCBR7rJDcWO5rw+tJo5Ten
NANhJ7nhaejaNYFGP66zSKmSKxyDXBlVocIxaPw8lIoNKRijjtb2I1hgipXL7XblB3J6H3lYoaZ8
obV+SSBy4xqrIHPVKMwRnnnMUqDo23ITiP1FgBFSxJ2VzTL2tZWTb5yCszNopjK+ljFRhZhEyGRG
boxHWuZIBNCtnLK56QcldwHT4KqCNnQ3AJvFP92TEuD0g8H+gNOd+sY3Vw3KBxofiuE8oKBfI0Py
GG0HH4UswcguTtXiPyAmKJ470GMY9gYDnvX9VrQcuhTocFWrXE98sCEvE6lQqdVqngcZNE7W7N7I
bfwqFyvxuTcv80o9aNEh4L0WlbaMX4WTht1bwrW8QlI+/+JlMjAge8Q/FBlhDHi/SfDPkE7WB4Sg
+I6Pm2w/oybdIb5ErbgTZubz3snkGGJvdD9FLGuTgQ8eKwosT9s1gDs7DKaGBaeV31p14mogTnaU
G5TMmUPOPxqahOWb8E4F8kFwHFKnyjC+4TQvlFi5Bazbjvw3T/UZf1ruMpet5pauC7spWvs4KPCc
00IJP3NevdIPzNo0nn91X8+OGelfwVSSblMmh2q/5v2MqAkV2oNWewUUbiQOp1OtuSvjXEoXH1Bj
HCjhHzJxferzKAKpUGIIuP6MyJk7unnzEsE5O2waPLEZ4YCztrUqIm07ItkBf1Bl+/uFik8XL87h
vr60DD9V+ICaUS5Xd8svWThuSk7BalvVct4J+aZskMgwUAc8t3LYOUfmwLzxvXJKeT3v36pS1QHv
OUtjJKiCAF4xyAOMyMUKwYeMhC3stfPG07GzGMweB4kCT1D5AB9+6PaDdfrZghA9QQ6RYexXuzk9
3Bc5esL5PJr4m/Yhz15ziBW9GbNTqKKkBmDMbaYshYP7eHToRTuxjtKL41lbioRLlijcFPL3Zs4G
4bDKUSjohhV2pPaK0YRSjS+Y86NnxJycww2Wyp/6GV0rzE271yBY1HA4M40u/pQDL3rC8KpMR8sc
pUG5wyS3HO5dIiwCDuCcOKMPGGqrzbEr+awvbkjBlDqH47a3AFNhR8+6rcaOdOizsIwYD1DFwqa2
oa8amuYnVoheKrGor6U+ccuJXamyM+gdEPGjvCGjTVxdAS9yi16G7P1h/xKVmitli7SmDLk3x9va
nT4Yk0U4DaAwp59MfU5Zl6ASs2ol53Ufo17QF6/BD59vOS3l1gM+jxsRg+Uk8xQ2c+jvXRDmpR35
NOTCFKy1or8ruhvVGFV6UITs8JBXY3NITBunQQa57u2p4xcu/tZx+a1lkaC/K3GQK93vXjdzYRIR
rFIvKOHpuAnBIf67KfimILjmR83PqwvPuSew6RSvssRqva9plER6R9V241j21hXNJKwJmrzmWWpD
Bw9qhw4wOvkwd5YFMIMby3WCBRvncPRRRyYnCObALhR5kmhZ8o4AUCm8aP8dstoF65uL3Jd8G3/7
Zz5Daf2Q/Q8155axC4Pl8Notz2AgaWpQHdQo3GLTwcbd3wJdeGzCyd6PoULiB9Uh432g2OeuP2Fp
Qtt7eZQCxVxPbRpvuNs+L5iEY5p6ItIFFQuaCdZigwaIk1C3lhlan1THDTSw6o0GL8egvS86NZZX
+R8Ft9EG40cJAz98vIA6tN+HZXxOO4iWoxfPNgEt3TR9aEC2Si9Kzc5DHAPvmhlKjhogrpNXIp3m
rAwb5Gd4aiA3JPMYPIHcyJc7m3ABsWgRGua3Q0eVDxfLKu0a7sMyxmp7edGLjulgM/xxd6VK/RNZ
gIKnalU77VjxV3okwVaPkTaaHJlqFhk12dijC62mZAteZEvQnj4ncvteiCikN7wdUIUaXvdAemks
jhENNVOfXfcyuuq2kYQgM0aIt3EeEtN2rP8yAtJ24lpJBiPy7r9e70hZu6gL6Le+S5yItzJijE69
h1HYMOzOJDxkdc1foc0FHFIgoN1Z0ws8fv77a5PGu1FDMG2DyWg29ZfMwk9prx7L1nsYR6FZB2wj
CElVcrlZBsG3U+qs3jsEKtBwsdvzvYG0MpsD2rUQYzSahWV4Yt6gCFCYEuZjX9sXsjkCDTvG1tC5
KTLdllAe7hnpsMsfN9i/8GPeQf1xgiHbdHoo0LDlbAtLs10BLwdb7bhU1o4Zyi3Ntio2/lsVvUoQ
OY3EEhk+vj7zEPjk6Q+jKojit3KWUmiztc8KF47QZWvLWJ31OOod/JFBGRRzVGa37vfkTlWyK+0A
LCEZkkxR1QvM6tdCh+EacgRXWiZ2h8Z+/QdpuU+q0LxoaxHjCfj/q9ILc3Px6XrrS8CqwpsdDTEb
+yn/ZQ8ThPd00GC/J3AREERxxi+6T9qGGZtorn5/tKHuPQsLei/rppEKLR5ij/aPOsft81uqt/aZ
6lqWDXCo9u49XiEAuPyk5H1o+rnf+HFG+S28dknXt8J2cwh49uoINjhmsMbFNST3y4eEHzBLctbU
sy6xhv7O5QPBkJ1Hz6eHekbX+sJ92NH5XnjyfRI0btwLCwjvJ0shwQWEPUG+CtSOrWZ6/ezBem9k
dtVba5DBft4hyx09DppahOloDHu7UDMOHPh5vdnkcf+o31Oj+y6Sqppp1Aj8YlhosBk+SIVu2NLP
qMs05nOkf3YfYdgAkmd14xnAJaH96r40shgd59MS9SeRd1VnTSI7eRUhhLXBp0U2BlCToGTjlhDD
LA/ST1AApvMSG0zbuNDYqCS2JEB3s9G1Pb9gvVUAgLmYb5bSvqNvzn0rklqVp5LtQVMjpL64/sEe
MgqYv0wEaxac9qilIJ0OMmyIbepJa+B9H/ZRcICV1rxOdi3alISXQzAYmChvPZzVd3R4EJ9XfaHt
/5x1Wq7ZN2guVyqHZ45qJt3j2cVP1KL0t6na23LsSN2twR0M7O/2Owr8goLiRf8dSC/Ee2OB1Yr7
bWLWQrGjumPTh5sGb2MNthQSowYkvNRAkvVKRbWblr7g3oi714yGVHGJmCNP0us5BTs7wbKogln/
UwFzorWye6y5BdQkEK8/p/5EsSZzPc94dIezdiL3nzMb5hslOds34tmDMDSUrE7f++HH8xobizL7
7gbjoTi3Iz2N0tXLWKjxKEWKvthcgsYWoh6qTIrsisRFvSb1XVgIHHCPkf6/SLDSn8x1vZGfNROZ
Xla+RNdimzBAClpAZP0Jluzm6Pg6QbW6oNZo9FipnMQmcXLUryG2mQVVR1d++BnMOo75aRk+CoB8
8D/RJ184jqZdvtC9iGshFvet7cCjid7GzbKPCvkfvY8d50jcDAflRWDpL5H/BOp8puZuRvDGmUYJ
GX79EAXhjf+NvO5xRv62Yn8hyzHhgXVIoYW7/2yc0F4xj4aCpImeGez0F5Po0guGxCGhp+Ns8RYY
NlJRpdeXM41EakfJYuZ0ht8BeDDsEKgPSYKGaI93SUcZV95pcS4aFr4MIXIDd8gi6fGrt1+mX62w
8vvcxecKRKBFdYWC+CVvpegx/QBrtoUIMfSrDCyqJwbIojsagE1C4DLX6rdZD5AUaW8kZTho/9n8
zg9FZbQDGyR/Y+PBJPO5brPVZalQIIkL9wZsH0r8gVnAZpSEte8GuaFEVjp7k+h/EQjvN5mcS0MU
MyKL1UvJ1VSNAVgPewYz13J3+uUKg2N4qgyBQhclztXhjwTyj2GeESohp5/9PCUp1d5w+B9GnJBB
OM7JsrjNPpNbiz+qfRxsBNAMcMSB0c9mtMtvQCPxeEJQgDQ9vwdBwrSJNn+zMS1kYGL4BEb/q+AW
Adu4zvBnVPwCBGPhF7R8WAKu4MQHN3OtLNNVwQyitLcQF7CvQBO3WsOBvQNqARMZc0CJNQKBpOXa
VALv7M2kat3WNW3sKYIi6yDxkxKg7zQOVj0CArS+hSVYvdTYb8LU5ZfZt9N2yEGEbI4zgFCD3OUm
xy6yMnGnaE0Gpa90vGd4T7HPvd/N/gCor/aENsygHK6my0XvfK6ODTmV2QCkjq5twBX8De3pbWo9
y/Uz2j5rE/YRoBxrcdlkefflT7FHLHzs/OsD3xSu/Evo+RLxIA+zP45xs6zhZIv1PM6eFt0NfuWB
Ts5juLdTsk4rwH6+vgpzLKiJVaDh2J9SzHi/FkJXtzPlA/ttOgKaWPgvrfc8cQr8gPIU6TGPeFIu
cKy4waYuGpUPJN0fYZQTe8B32lXPGmaMP7seTU5Jj/SYbyKMVHzs+7/ZhMrXkzkOAdj6frijYw3m
HU6YOWOPtBkO9qoOmivacRRahvkrIFiUwsXdqbDiCKhvprT+qubgYjUIb1xpN2l00Mppeby/y3H8
e3plcuraInnN3xbXwehTGJlmAQMX5HdW6LeDzSPt5ykLVg/f32MPSZcFpNOa22SZu8Z2F1zEZjpD
e8yZe9oWfZsuKA50gfu8daSfmjTKktTJZr9LEfslVRs6Q2YZDq9LWKffEt/OdtIZhXn7CG1wbECe
codDBaQbDRrj53RUr+1pq8zok8Y8ajfLmf1FZjxBU/rs/856jVusbEc68Z3Fw5VI2aIu0WqM1koc
6CyZLS3Y8Axc4du8A1tLsK3CBcwBdm5dEA260hr+gaq/TPnilu2WHqpR3t6wf4ZxFiEL3SEMIFko
z0/8yx2s9EBOMLadlCr769dI81EWC8Uynooj/q9FOuunsg4Tzlss3zo4JZJlZE6Dwae5PTR/4NA4
WJDGA8T1G2jEMXY2ELgoTbzrKn9pPdyxREJOfwVSSFVCGs5LVySaK/9Cpn0qDdmTKbALqUlic6YW
ty6Rr7MmWeG8OY+2DD2Ja6FJe3ORn3kj21/IFF0xoFT+IbKH6aJ1zO1h1DCceFSq+PGVFnvF+wLN
u+g5tMhpSowncrtfLgXRCbaxgn6dJIAoqSyJozTJb1EarIQYLloAtOrHBesKuMRIq5i5a/KMbTNs
KrhFSQIYHKYu5zjKlipcRTgkbIpmn61l5G11/CyNJTXSceByn6cpd6bGIHEqkxNIngHyFNPtUz6t
Bf+56IcmcvpRJ8fcDbtudzJN/XMMI8l4APTxLfba4FKYQNQJlWoLqXTMZzRTdGK1axHPIoQ5UL3x
LuzQLjOoEjok49SR64/Ivi33MASLCsvAZBvG5puSs4e5+PQFrhgaAbqrImvc0vMXrjcUagBm/xtB
wSyTFla7Tt0KqCjF8bk2rYaX5ayy7XUwY+Qbvf088alIPUrBJ6UncR0iloBoSP2qvrnKx3pZfLT9
eWCZdqpbCqyF8tHyELlfof+E5gc0u9U79jKE861o8I1EUpxFWTWplTO3J9ZvGDxRemNq/wseALLv
1t2xDImr65blRTg6Hw9BWEtFgmy+I0niXGTyuFe4aCWMUJB+6fp3U64/jrnfVDDinxEMNiS2B3Rn
jY9joFbXU/mn82KaxcGm4xLo3fXEO5nYm+Tfa7cAbmdlDt/WW5NRihN8rDtQwf3dFXMgx32EhNyu
w/rSMcRjd2M75QjF1hDXIwBke1pRriku1OK0cmVhfccpolaQWvWtqO1ZPdKbiTFgF2u6JW9yoVCn
7AuxAdyvxLIG1Lr2sF4yEccJa/rBVL/XQtJ5tBaclm5D9yEiNy8vhvjnjzk/oPtdZOkc2YMgsL+m
fuMGabnZz7/BiGqWlot4ff2iWGVPB+B9Bsak5/aRvUajaxNZ17wN4hRyDTAkRhmDUGgn9PDWPUN1
uzD53bMozBGOXICcO+iL9Fnc1u66dEoepr0l/GvcuDRmyYvqMLZeadTOeW0vzMgWpaU2fD64Qkll
hxA6BLb3lUjso4OQEDankQX+TqqsvXwNqU5DX4NishHA9kR0fRTfqGgs4OB3Fup72H1ZaexX7+ie
3RDqp61AyTm1G55YSoIx3uvUHJak77+tH6atO5TTT3+ikD+Y5DcYxamoNtYfQZoI7AOnFEZaW3SW
IO9X+tE9IArnZ0cKoUqYMzwXgYpMZNU6o5ZYSbWGdmpt5mnv8ImVhbBkU+dzTneNILnX6/cph9y2
ZgS1GWDhl5qRdjW8yNoEHt7fFHppye9hGiysJjRABpdc46wHZBv9ZAh4NaGu7RBYoIQv2EWEPBs1
qg+5VyCfrjmhQhoKXsScuPFpvPs348qD8oubygMP22uFPaJdT73p3/Tsr2xyyebNfVJAOg3g3FYS
ILs4sdphnnNfgK80iLHXteM5Y5AgyVjujKuGHH+cdYoztPDKE5+7CQBvX9rmQWdsovx/WDGRJpdf
cQ5WNHROEX0+BpiaK8FGXcyl9vRqeD1ndGcZm97F6HVrdrxoNtbeGNU6FAbTs2m7/QNOSNwAcaVz
vpXVGbjy9pkBpbss74F2po4vNU6jVvANz2K9JioJY97BSi9YU5ryWLkrs7tyawKnEbR8yYeit2gQ
FHS5b8jbkoQw0nBPNnmHnfh7EFsnYY2RiHeieqfd1RIzKN05Ic/HhTwFaVoRQ+4Nm1rwv3xeT4jr
4b7DfpetktU8brsImCKiR9L9/VdgT3EY/8UFJdPOT/B5bqxjiMoDSQallJOJqjCFxs+sX5Dz40s/
htF/7uhiUnC82pzH7WH8dHfJHBRnWP0IEzTe/jgyKCZzCUWRp+0lXr20ZpOTcmImH6XmaS2jParb
jkqBesCPnxBVUOt/BzgbOeXUSBDEMfnm7X1qyzZ/rPiSpmLfjZbzwgHOVm5LCmjriFwvwhyZe4hk
/FSgSZZqAGPYD2BGcoOuOv/P30zGBVYkxjArMaMfC1GSHCvj4a652fYdOrm63v7tu1BkG0bGB2w5
Ftb9olPOnifrDYsQ/k4ogtFkBlPKnPJKhGe8Q1UtCMiolalGlLdEmEIDzeco9IsjARrj+kTQSKs9
KS5oEVSxHQhyDc0GQ/27vsWrZciN3CVZeFopqqyAyHwb23VXjTkCKrE6fhFw4QlfQflX0QwGb9hz
CFnMfahbqjfwO8C8yxULEeZamT/g+P2Dbyi2NRWaLWUZiMeFAQRHLKT1aX7uD/tjbMBuFY1SKuS6
b7Jjb42h6eBeJ8S6CC/vO6bKopbqSSMkG+9cY7GAOorRIxMm5agBXq5A66rJrF8UbAYQ3inTOWx8
ECepZHWp1hQeYrLH4oJiFsAQNNn65kVzKzprDgL6KC2zvoiH/go0liXCpXEEYtrtv6/rzyvmdGqU
fEtTBmGV7P5fI4iaRlCTSVY/50cAEHWa8a9QPZk76YVCDPFb17pyPwynUyRH2cVXMvmOXWqPwWUA
TOVsc8CJ/6OOgRgwaR97+A5LchoUvf78usOQeHY3i7FmEbozT6IsqCPDhIpegVBV3Z04o+heft+x
GHl0WSRKEHsy69+RfXoTnhLYgrm3pMoBqcuaJKAojpcb/Wr3g9G6GFyYn3uDiFSqKjN4xSGuZJXr
JXuGrH9NaAoXghKuqZ+N3vU1+9RXomuKmeIxktOnZoM3QpXEZ489dTHzf9gcOrWQmu/mkAiknhhu
21RY5fdfVclMbVdR1W2aVajs/BmuoWdipcRRM2rV5hejbNMTmsE7BWvPOBkFYk5eh00teOuojx7R
d1vY0Lw2Twr3VNjlrzntdExmAy+02Bd04Nxe1RQUZbxbGuDECRA1dTga5oemCViQuXtd0A/kPp1G
zRZOGPkyZpXwUoh2PZNkh9aBpXTTlhUOq3B5h6Ke4Ljg8NUNZhfmh1jSXVq4M4ISpq6jSY/tHNa9
mp3Pe0HTgznMQoJMbKrAH/RaLKO01/5/LYn8NW6SZJdorPUpXIfgBJ8NvJ5TVC44uKAbU+f4Jrav
Ypd74Pqt2jOB+Cud9dDdR7kLTd7aZ4MMy4imI5ZG7zktVYs3lA6hzU+DDys83fZydsiSqBAYn97m
rr/YoAUV4gd+ydq9ciUu6IXTmv/v171Hxw3OBr40wec1kwfsmWBmEITMh3O0mZsX/UqraWmjB2L/
UzWQTtN/emSgZt59Bx5CBAHgFYH5c9MOt7HbSHY2Xf6fq/3HVTpWtDNhL2mwCEJ54V48CNpypcCn
snBDPAlmbGEkN34LObk8fkxyibBpAOA6nG7wVz+QvpH+ehiKQNQwaTZd/zF2OcAanGpVNS4GcKib
wXTuPAIs3rxEkATF9DBg50oAerJBCVqKTP0sJyrblDQJWR0a+eZnodlRlndwySFslvSy1gEARn2N
DkN4bidmG3ByJzAFpRoifITYxrIRw9WU2lkDN126iyAwEboEcLfms9KgHk4cgvyEq1BXO1pYsFjQ
/La1YISKNgx+xiPQYY2BQkspgDFCPlWwvKkXsSL9hzDXA6vBNs+CF49h6+HnhoBqz8JeRbrCWhSj
Ai6pzu2afBL4JMNYuprNdWUvd/XO6HMagqwbNXIPLH5uldc4BYJweCBeVQmMA93upiOcEL+wUB0/
3NT6KKEioaAsGCg5fMPEjLv2+/xXKf8s58B7Pc9PfBe39CYD7HCCt4vbX5HzRaq2GHUuHZ8AY6TQ
jsuKwX69h2mXE7jRUZ68aHrPQSPsKy6zJfDfaGmgqxCpiKFIXzwx67cSRfk5HFu1GRpjcaVaR4p6
JoKHiQaqVRIObif7cMIDaX1rG8jaQs3nFalJoskLRiByDZC2CNaRCMVyHejhLc0Nb3sdwrUDBmWe
zNjBiBE5GRg4Abxi+yVas8TyOf438dZTWmUGfKUL6UKBnb5hEcK7O/myRw1ScyW9xju3vDxNwFMu
AwxoudW8CxzJHSn8oCp1v46GNq9dzTdQrkDafL2AuzYYZII8uUGVisLeYG8pZlCf7vDP+PfWYZGy
33c43F6P/wwro0Uw9tP8EP4rrQD0EcYpKo8W9CFjUN+0ylnYsZTCOI01j7cXTD+JQI4qIVW9w1mY
ILt4+MjeL4J9vj3727UnwYN14Vxdd71nm665cwnzf+Q6tOYXbFHJ6tQi9IGE55NwUNogVALI33np
jTKfk24ly0M/DtLvz5cGW30u6elVRVPYsbwCJsLvy60pJe4xY14OFEl9qMro80ppnQIEh7hos58D
UJsjqdE7NwEMNxyJHLewSVWBnfZWW9D75xLDuxKHsFTMDbl+B9Jd8n5CLQcn1pZI83JccJ0UJIqc
sOu5mcIVwuZxEXpxqvv/01jOdBwZybaxUg0Ab4v31eSxpZ4ojba7EQshEAYd5tWtJS98FvIIosE1
z7Q+s6ppRPYi6ErizjC9iOZpNJPW+NZhrfCQ9iSodMUqgd5pao/IfKIaJGBz9krYk9ZP+h8dVC2l
RGVAp+hNGXxvp54uoKh8pjAaMS3XqASrveyLjwILOVbGH7fzr6bAU2Ntf+6qrLapb/q/cMQk8g9r
yPil837FqL9BkFtu0L0upPI0Bm9bh2Wn30UXapl36+VIzw/o8r243G7MdKVMn2NDP0nHB+TrhMwT
muI7wlMsINevQxKwCGFHuNk7rYpiFilVnyzz+8IiFmTNwZ2dfaRa03xdEbdzKJji/JWC9PPVUMqO
MvDlNkDSb7dwyBp3Ck0FqO6vYi2dT6FBxmiJq4AAoNzzoICjZcerD3GF7Qvm2zByWfSosFdV6+NE
liU373s93yjUQvKavP137R13wPGn64fI+pgIvCOYgplztA4lTecZsrsZhjuoEFxcsm7FZ1kiswrb
ZbrdDBgloUpOCVdjJbqS/pLY5TzwxaOZ0MoeunEI4dMbHB6t/aC3+dNvQ4T811OjLK4y8b43pbZZ
0XzRcZdKfbDU8esRb+X108dAj/3eCBsOfCvV94c/TGJ7DJnHaQEL1LYcRr2gkvTEhtiAfISuxgMy
8OukPEtHhk6JGY/ZZv77eIdcDaGc0yfINYq1hQJpTrrRDxaiel00xGzji/e9eZaq2oyEKT8uD04Y
A1zZqKvFzo9ucWamVFFX/vgs1nF2kNsdjGBhxL+9bdJrSCzH5fH1La0diJpf+rh8Cky5dkRsW6XC
igceb1BzAIPElSkX2YvJ/ElWKRMvBslBaLsbcY9whoIQ3CGfjRSjMrnYFKYUlEwu6H2nUc0XGWqU
IvAXTvjquYbHAsiA8WPNntQNCnHAHyP8iyuXnchzsHUw2PnHh37uUgoVn7/+iHl4PnfHbkYRJBKy
UruetmhwW1QIRO3k0TZF8UbfR5DtBoO+X32/ePVy2sdJsqUHsWdSRsxbMlrPCTGYAfNOauFFr15/
Yuyh/UlfnBiXg7YhRskpkwgfvSdl6imDyGImD7zdl95kd3ZuDJVBknSIfC67q6gqHEvnR5ObdOew
pSK0Nfm6YX4/cpTydeFFBLbGDIH++T3wIgvueMEiVBqhEjeekgqEDWTohpJDiyRhfkL2Fu6SaA0g
2mQknmrLcXspeRAeo3tRMqy7VkWgYJNf0fSpz9pPIN8CqwkwgRgD/2GP4MM7Q4uBfSktDrrqmX+I
0aejB4k0qxEDgJjpEV3s/7OIktEGVR2FjtlhmORwim+NYy9DvKrCLNuiqZCtD77QXOY8nGRXlNbs
MTXm3RpeaHIenSWYzYKTVuhFLuzxmUTY/JGkk0EikM80TiXs+O7WXmNm6bO2lUjn55REowN4gjIk
px+lK/UL7vhJy+aSmB9kvrpNHeIe0hN0bjIMtwb/1HUceU2LpQf6s29Q4ZbtPDZpL2jbJ2vvDLd9
Nhc1KBnLTd4kY6kfmQVfJndrS/oAnt5vky+H3nRsr8/oFcx9EaLf+qEdeHP5RKa1EiCu3qnfW1Lt
9xCu9BrfYr8QJg4/RRQByxhUpwP+ApgPOO4cBDbcTBqdE+X4/u09gD+hx+fMHv7q0WNxENERt3O0
Ydq0VvpWZIU3pwYJVQ2rDV345A1tzOOySuv/dUDoA8qwpBPeInW+GhT5PlsYXWf9ezCATSCUIzoJ
E/QqV6ssGdv6V0mE6uqDvDxEpAlrvljnSiuXF0P56LwpmlkRgkjYr5i9ZVEFheACUDm59Oadd+Hq
3wsHFF7Gb9lay4tYgA4046Cy4ZmZLNWgOccWKJCf3djSon2VyYZPKgaJ77uGp0um4jloqeor8cvS
0aTXamyaRYK3GTFiAB25I2YnmaD74Gp2M6+hxvST9/V634wZbY3156r2rfQGK4pI40pOS4eRYNf/
lN7Gl6AmYm/537+pp0k8bj6LucnJEuCZgaj8wPE4l16y0GqNMiRWSLFDi6FaXftla/R8B//A7kEl
iEipNcOY9vGxRtgSmeijati8RFsDxT9nH6vtbOc4mYOsPX6r+aeUxnL8RfB1n/csSFQAdrbzSl2P
oYN/Fym+F8ZRd7n+TEcHkY9awd3hPCH3ZHPLGCXSn+iMQxrGay1Pdqdjc2p/2F2zGnWod3BkRpU4
0Ldl7Pt/Ryc3xmkFKaQU8T+ySF9yrDV6c9DyR1FKzxvxFd60gw3HhZAeyDbc94+n8SDIOJVh00A3
1QV3Dh09txBnPzJ1FBSPuF7al2fOtFaYFHT2AYhu94XWJnnqwkbmt0V2RPaA7sLkM0YSQXM89bUo
W4gaw6oGDeyHuT6LeBX0Q1+TW1ABB7ktiReWYNo0pG5I9vM5NWpixdoALvLNNVkxUZYEw3R281Go
pkF5OjAzejWnLOyNxXZG21b4y6ssCph89YKOJkvMDjiLfHUepizowyPtYEssh7wcrd/drYnsA+1m
mAER+pfyi6O4qOcleGNDAIXyzU3JROiyfyZmwk3f8EG/fjjqR+DDxA9Go43ZWNrckzJIGG5/vEYz
TiMlu0/wGJMtFA3gSKHAluTgtGtlx/qKDWXZzlI7Lzk4jzL8o38wwWVAhsqgXgr0LhpjVSQFKtVK
qL1JwPaHuqG/JjECg/48Jb6Dl0C4GTF369hykMGmCKicfjjehKzpwHY35YcMdfylvQrC2d0P3IGF
5JIyjCPjlPpbnihwldKO0WV1Ugj1CTnZJ4Nun4jbTpJhGHJQ02vRqnqf0zPkq9zTgiKyp7PK7dsQ
gTE7zTpg8+zLW2qJ57klmUQsZE2NWYXLMyxVEXj2I4qm+pl3CyTIKevbz4EH86AxfQ9D50TdSEzq
aNdE3bdfef5d+64unUyNRjqIMb0HIlptjI52mNm10ggXo9zQtI/Ner8aKvIvb256g2mtgWlTdfGL
e0bjEK5e6upNygunskZqzimAUf8OJRcEGdGNFV0hlwlkJ9E/xrj9/WUuKK4fvNW8WyQk+E5Hj2li
680rCCcchvIxChQQaFrkDG1XEv7nMNDBjsgZxa10RvcVrhF/QroJHQSTZLcw6TDhSMe8iW2fD0Z4
AexZHSmovs6ZGt2XcbnFNo+aUToeQmOzeDsU7xlJajZueQ/Ss/ns2ExiqwwXc2VJtoPPFKFcDYK/
9yao7UuVWKLoJsxfAVO+6H9mhX0mBcoQqBH9q3INfZiBq1aKl0CfzvRwhQGsRwQh0nEKEnDqOOmD
zdEjiUdO9d6RSqc1KXpkoLRpx+pk44EXG7La2A9EGOjysHlWZTULC6uTukSgDO1JXfHWyCb+rCtQ
IrmsMjBVSWok8nZpbP0TLtNVoO8hAgMuwnqKz0OO5lb4M0MQfc1rZnupzq+UhsyRnX7iXjTNMa/6
RoELtwrHLk4ThwLIOSOcXRE4dXXZQaDK1oAvmOyVIyxffVo3hMOiW2dyVUIsp5ZaWmtJMsjsnjmT
dbLwPL7jIXQjn9PLIlimaQZf3pWE5+LvYGUgDoScofQBQqWsmL6ni5AK8+SyXuRtX4ZPYQnqgMzC
R8fQ7kLTSyHbaf2bCGbh5TbFrwzAO6CNWb4cRU/oBEocSAqzPScshhU+JrNajPSRpWYnnvXe4JlE
OoyXVnIVY94r+Cp5q6ffrIYF16XJRn4GfxpikF4mwGng73y+0w1th1/WjnH92b4zPtfdgeDkbw/8
99Eo4402dWr1DP/YoxDUTPNYgBZgxZvIM0g4CKlg5FnS5KVLT/l+hPoqZa/tPuw55w52b2WdOeIU
ZDQuhy+w8jrbptPt+4VA4SRO+I8h7y5/rwfeO3EIa2ZUowNi14bQ0smGUTo0utlG85TZp2whsP2Y
DzMrciDMSbjnx31KWKm60Jj6z+AnrPk0hXJhVbVFGmXCRZA3EDmVP80INsO+ky54wUflxIsPkAZ1
PuS0u4bb8/fi6TRpFJyrCyKMeEwvzC8V9roySkkBwatr40ChidetlsFY05fe9FTAyQZjz54NmakA
EvfeReKDPP5ompR8SWcWx2NA3SaM1tAtf4cQ7I+OPPo4fOvFN3N9DKhI0Mb7mz/N2HkDWjb69Hho
+LmAAU4PkvuUZSIHbSDhoP/QT69XDuUfL96P8A8SCYj7FeWEVWn26F7DE55rTBjT/iXtm4GDRLu3
QRHWnjRF0IB9t4QAbo7G0+XPM3CHd8LvdyTQOeDav7QSde7IrOmxkqaAIm5Nx+48iL/DTrEPcDyW
vFEZZOt85B+lMtkLYK96CM3+BgLUqwTGeL7SISOptC0xztpMgqxeiIVRunRZrAdgZrSjacCbHYGz
c0gWr0cbyoeJqyFRnNzJM6xbdkBgOoRmavEjXm34nOZnFGWdvbLT3U1ZhZPzx7KqHLKxs6c0k9HA
tfUDgSAQ4M2MJ/cCaKNf9ZIsxwYwg/7antaYQdmKsOuJpOPaS5Pi8qp7mTnk8DLKycEEtVU/pxXv
dE2oSL2UMe+GgRAhWQpkDqRdbzeLVUayDagsEc2bcASwqj8ZvNVwYZAgzY1/wYryfEq4vTgAaomf
ik0PXHizBsNrE9pa/hrnYQXZI6Vn5KHw4ORwazdBaeRbC01hEMov1zBdnYPLRLnPpffs4WlqE0rr
dgx+GYBAifhpyHBmfr9ajj2zwXD50zzyqYUpTXmPQlW9Py5c2Kji4p7fx6wkPDXjVisdB/c/noTa
3T76w5/ppOB93RkXqU2ObSX35ZPg966pyVmDRMb6AIP6o0lhlr/SYIlD2Causgxdz+VfWvp57g58
Ih5/H1tS9HSV/tTlkeo7x1bNF4YDvAeHVspyJ4JG/3rbPHIR4IO0oNTGQbQUGbLL6Yon6jjhdJUl
NVwtqr7fdGKglng9bbAOkO2T7yMOQxTEYSyHvJH2BBmlKC6FV6nWx0CXUon5INTrwMheKbrVTBZE
WTYVnGqLUWS8RrnH0Yaj06HgXCjfP80c4YjMVMg1jju693KxykdCJHUyLzGNSU7nkUK+U0S6PGJ9
K+gEJ3A1D7Ywi6iDJKM+qvh3WtGAeerMRwSBPU4i/T6kPT8ngAovH1kAXA0RUYkhwonfgV3NwE8A
DmxMGucJTfcyphVVNyr4LaxmDZAKvjfKi8NShKAJ5on0rIPbv/Hgz6bd05etD2di66jWqataHiAd
jjIWjTLti3pe+Jfa7pO453SeVJvj0xME1wGQESfrZVaVrUlzdWRtdqb5x9HjTcPkX/lsHn8eMoed
HKfvQ62uorOBqGATLkhFCp/QOxvEeEatqeliIaJDLsBRzW4K/t3k8D7tod2Xbdb7Vv8Yv7BUQ57h
OAym6OgJKDHoHiUqJiHsoqRFal9wbBdMMEJfEeoC1f9wkf1Nj21Ve9VtA0RigjWL6nme8wuquqdM
bgORmQAOGUxW2Eon4zkAURBjpjHEYhl9I+K8uPvJUkLTeQZEj5WU/arM/Ces0jTBnsWrbVJagdQE
pN/drpoyIJ7rN5ksJXAXOfXffdb1rg8hbBdSBpVeMfSxwWR0BOkPHD7RJv+X7Zy9em7tZtYPHuAD
u1mZUvpiQhVQrfYIBVR59eYy+kG9c/tpVAFJZXZvM6eGivoF9D/HqlHUOmg5t16yvY0B+j+GzFhx
x/2fV9JZ9oTdk1QkKhpOHqISCdhvVaCnZA/QemQ/0IeBLBAjV7xLcIOJKXuEN23Xt1d3nWnMdVkB
/Q8PtDfoZ3kTx1cIfllr48bMSOvYbR5xJ+UqjgxhkXtSj2S4UsxPjx8hXXFOUq3SKwLblpucj5E+
kSool4POpOpZl2K30OpkcK3NzT+miwp0cHCJ6+zcCLG/nI28v7LgUmtQXJlm7PKBl5feLfeiowyu
4XsHbtl8MOhR731RmB3B1IcLcL/XqQ/nfYHxdviiqbWIUBuPEozDZP1l0gr50+4huprpOtfU34Ae
aEI1FuFydaAhMpiYevMW6Hh91CAaJL8z1/PSDX/P2VDl5SB2Jnxuc9vb8EoE2se3y9yr5nVHzNRt
3a4o5Yk5zAbJbSKu6iWifPTsRKKm1cvicr++PSw2ClB1PuDZUVYSCRbqpz1D0mltkoIEkO887Roz
HnPEkA2VOMd7eBf1lEbIDJjLM8XnHr/UA4yIFS8JlHokLX7Mew8AoBmIJtEvXjfhyjbxe0s/0xTs
+BvnuRF23ZfpkCCikuF+yDQFfPZzakuNT98LHzNZafzJ8FKgClXaZUaPH4krIqWKhi+1PT+B9TyV
6qypRfJQo0gqMdwZTg8ocNzgY94GFoqc5ADgo17W2tuvaysdSUdqqZjrsQKbO2k2jiDKG/fPnnsu
39AgRy+Glz1Ox9WzPC89ejKCBx3ktCeWMllOnvl4Bzp0rl4Nx2bMVc0YhUMYowMT01VJDz5R1xTa
dTJ1vaKSY6iXgnFEO3GNs2273T/Y3HHeNUgQ2QAlq7iUDfwpZGS+sUBM5GX7RYjCpQv8u1tVNWDC
rfGTVqOD19XpIzrahPW5PDvByxtEyyjzGwPOKYWTvaj0pjGFk+RpXvIxSKdDDJnG8nycl6lAZOTS
3sLPgSVKrZXqvYINyWAIaoX6MFQx44phEXYibXJO0TXUAMKSZvmMLzc5A3+Q8O6vH38f6J9RC9cL
leleS0T85c+jcKSLWlHHpEv7lv4UqQKGIWahzYeN3Vw6dcCcnvFij1l2OUtzHJxq09jLg4Ia8ZMY
s3XB0yHM8TNTeHpqMNGgNH+G8kOstEeMVZC8rFR+2PfRsJnGDVYBFQMdAwNkRI5q+QLarTKaZDOT
UIR2zUW+Wn5R86+nKqsviWKyGR/W5Tm8DlsR/kuZ0UUfaBYy8vgFXp/sVY4odaaC16mPbd640ZW6
QKC0y3afNZSJ2S6hYCo8dOHSv9dE/rw1SlYbf6DavLLOAdZBdTcLSss+GmCD8vFuT2ABRYlwZiUO
rXduBBi0CAwcXR7c+XN85G3ekls8cXtF8iIXrR7CvPU47lEaje3G8wbgrYPLPf7MH6nnZs1Xv/rr
rbyR3RBfZ0WjAo793xNBRcnx+ta/8Da75oLf8iYdmiMX5mQghgwq8qTHoFgXjRRscHn04v6V5az/
yl1tUqkkvT6tiu/dat2QFseqv/Igl5ESjUSAXUN5n75Q1+EDymY8f//cy5kAVZ0QLFmozOV751LN
gFcWhwlunPUwF7xX3N8EVyd8WEm7MBnxwwZ7USux4KBAm1fGHROUNpozzuZbg0Y+zsBFzA9xWLGI
Pf/PUNxoDzo8YHsNWUEXnmOMOyJXSvEav5XAxejsJvA63N6eDZJY/gDVzdJKVHTfxaAG8wnzVe2Y
cblrAdZgY7ZTKWAGS7hCr8TJVhKMP6lC52ans7CY2jBavRZw0+TIyISvYTwVMY4rQvja8MnefhYe
p5C3G0KttaeBvSH+WDapibPMe/EHFW+8b7Y5nNXMnGiOQSsEG9XpYkgdE4EegYAvD/igIpYzy3tI
a7jyt+PZuASvoweoB8GVPps0jbyGy86Xnc9SO9LcbhYAKil+uzqn8JKXsMxR1Xbjw6rgxYjGpwNR
sVKjkm2iHkMh8RMIPs/h5HBrcS4bN68GWnje92GiDtgAUazSxdIAJ5+szC1d8V4w6irDMY0jLyHn
2b5OS/GCj8RoWi7ymZIHTXJB3+lIbKQk0LRwg7YWRWNpbZw+PC/udGieD+G/DPcYrbQmeV4gHWwr
jyqq+6c/+qrFTywD2bcgGuvLbyUpTeR57wKCfsUN2d4zodZdfekgtmdzt46afaP3fdyHfIL71Uu6
py/kTrbLqUZmrBltBhMK4J3BMTMmyD0Y75DjiIO5GCmVpG+EY4pzYCl77lxCWP5YsWZekEvWoClj
J3LUUe9Pl8EnwrFmySFbv2PpIesuT1L9o8LpqD1pAOCXq5lAKcwSrt9FVjo7serhJP7E+tgphKf7
StgCAJYLPobvWGcjS65XlJWfEUE0c9xwy4s3eDOkYb+TR8UdXiBE5B+zunxeg8G2px1ZV8/pwmcd
MfYddNXeDCoovRwfmGXpCtzN9dRDwKkvE3gUsE/QMBktvbkSgboFLYgiGOVz9qhNMiWgBSR/vNT3
nG0ZLaS2yVRhNIWmA12fPBRIFEDQjPcsEEE1Bz1Q029ITMc/OMWVw+8e0vTG+RJoQ1jOfgbnj99D
7TAo9gPqxvpQ7cd8y8bdnUViM6dy+KeibotIAg3ghmPl4QfvrmjBjAF8Vk6vjE6Nw+HM6D+s2f/I
j/+tUSi4rnCikyXKWUJZWyFQ9LBAzsDUNXv0iozvPYWpSgvuYshNxF1IqG+KKGzSrT3I8qGER9XZ
LdYh82Fc8oAt6Z+YVZQ1pmMNLmKD0GajGVxFHWmdMBtorv/8fvft4hzH4dgLMndK8UEMnD6BT1ZQ
z06HOnYz58ChBU8zlAjn1P89B9fBqTWCEnMG4r8gZWcgtIxbYiuif+FHI+Jf2M/RseYYhrw/rQSV
S7/t7yrkL05MyqU2lYGSxOw+Kski0oZyJCShwbMFsdsVnJb/nm+OI9u5tzve0HeSGVL2PK/zSQC5
X0urlFQHat613V5OZPVk7ZWxdUzUjfsB2AUUnNKOepo8Y3SPbitiK/vsCJ8J/E80vxEHRN6fZvEZ
nzM0Lh8HQRh0svS5+sGUcpuJtFIYQXmCLkUelhEj9LenvpkYm/0LzKNzyIMK7bVhlzahaIKX7Pdn
Wz9OTWC7J2AX/9Wtm8vzYKFKgDJg3FOOFtJDDkcQz+f9z7rz64u9V9RRQqjbobd4UYpApBp9Y4sv
3Kawj0IflVtcoGidz3QyXnqS/Ii0rwCKxujnttngIOr/lIE/KVqDCT4+Q+U94OmFXjdoWcdPhBDs
2lSX+caAS6MLvYt8AZCdTFuFc/HH02JF2lVVSakb13w72Yl2Wcw8lcc7rMgOojaVOxMTSqP4oMl9
e4wvZDTJBjK6NqNDK6UjgUbmfSbGgmdIamSnpBUtHBFlClJm3hW2A8dGvc8j1NrFnzDeMK9NK3uE
Qp5fzcB3dM72lV9UQLEtz8Cfi27TmtbdEmQEtXL0zTKlIHwUvMwcZDziUPxcxvqlIH4DrMfSazz/
6nmtzSe8eesFWFWoqHPno0L9L+1sPMYARSnyH3ey1Yea2Bxc+U3pKSS5EtaR0TIGXP7vn5aulXmQ
5LhS79wXAS5/PXdETkRKNWVIDVVYkElx/tf7+WwFXXSqwaF4w6QIHaAWbQtLbl51QcmnDCeVhI0Y
p93tB/HZFcfxnHZD/rm1ChHrtjXGTAtGMH6CgRnZa7rEJzG9jq74kPky2QF1PRG3P4rn0c8dbiU9
JTe+9brOlMS8EBZjX+smR6XTW3AFHdpFXk0I442skOUaFafMJaZ2Kb3PZG2PQsXg+emmq97NVBQa
pg2RXXF45mxS04KLMIlJe1cVtTFP2IEL6gfqZEkqebKmL4ZNGp+2cOh3uViJv0SZMS7T/xTcfkhc
SMlGTJMebuLyiZyfa/Ju6sCgaWKTa760epiTzuU/NP6CdLrS//s5BNkpvWsHAa9PD15YgTYQZyVq
gKYPy8qPRLNdoSLS4vYG15lAi5LBEQ5qG9kLE/M9HHMcrU2cZOccwg6zRwgpbQHMBAn9gr4Hegk+
5y+qDLv6fSCEAq6Y+tgfoBtuAcIyTmVAxztstbVoxSCssZ53lbD1BWTDvKooD6C9LKIXiL3daMxx
IX0WZlWTbk1fAqcXUyZAB+bDPlGCHMnH4eXJyhavx82azrQOuC6VZGG/I3hOvch1fEfxgmBsq2T7
KK0Ax3TBBvM2AWad3Vq2Bo1dgVtvB60rscNRpeBTqFUcAW7Zq2z0f9gNRd28Pf6q7Fk9VNLXOwCN
teUP/mg+tU2Af5D3xyF2EPBB3/mAI/aZY8vaRf4mP1CdIzZceuLX7NAT9qkjJS/waJfpDKkjkCyn
Ps0m+oQELnuvX6E06q1egYPHZiKxT7OO/ea/+yEMQSeddHGqvgmSwBHFodlEWO1fwOob+ty+wWXk
/OLfKaU2HMHUeicBeHhqCoHY4Fhk9ISluARNAjHDr25WZi6YJ2AihXEb2juR0EmHjtFZ+KjeaeZr
Q8+LnCKyYrVJNWvZAcHlaq67zt6k3MHiGeD//fYeZPWjFG9LncHAeLpy4qQ+jDOdn/zGAN3GD0JJ
uT//6O3c4JfvHaeXUR1djVN/cLjrEw1+7B35w7fte3y4Y/QMXzPXZteYc7iNp+28P/7+xzMX4Q6/
qT6cujkU9FRuYpKl+/B8gRk8kjy9ZcdKyzU5MfJcKSzU3z0SqwiU1rJB3+SPmIyzUufK9Z3Jk82p
JnHoTskvQe2r5Wr5L5F/SMI+K0eZ2tXWVdJnoyXsU4P3oa8VlrTM8QRwt8NLVWmOm+2Qy6JQQjJG
kH6SUPYFcRwqs4MjR4kG6oQnwGjxuqQa7Dfb9IovWNlxbAlFrv8U1DOvDd/qGZRt4pHzpdYjO4W7
1B/sHIOlbiACzguKi3iar0rNQAy0Db650Xh4NpAohbFKU8FnHrC5tX+pG4g8L0AUuvdSwzbwej1N
r7gt3yCNj/RRjxSxlRlym0kxUhsNeuiRK8smYzV4KVeIJQzDAiHvlSwpToFjIx9pCfmxaYdN6MBF
dh0EVwMoxKiLIcYNhfC+Iir1ms7vOR54kKQMX193q0XHDo/qoTZCTXmSumeXcqEm2JUN9DsfVSpM
Rem5FpNU2HDyl/TpI4h+ElFn/GgSwzp5KK9VqyN5yOA9Y7/CyRr1K3uw91UIDA7T7gDyqQhRpI9z
HNMp153nM6FRWP3NT3TKkJUXxmpTjNe0ktFqMi2tAPRkUMSeb6FdPhVdwW+nndEaO1NN4dEa87Qf
GHsw6RPEYkpD1gMT2iDlTIe07yy6Vfuf3EZtKof3voPD34Q4kJFvkC1lMnViXf7vt21866lU280s
PBKwJwDP0jd5tu3Rj6iqrNSvffb1XZBrVRsUDzT7VjlM1eNIEmnLYDAI2wZ8/XGWmJI8nSi9bOp/
EbfSoOny3gx9MAjfcJuoWLkOnLQnEBqrGzjFWKcgM4MSMIzcVRULyVhAb1nNe36GdWg5dlSNmT6g
ZRaKt2VClSIBVMnP3eSsL+szXKZPm2PPKA2lJwrrfqQg5lbMt84z5tcpaXkgq7lnuwnsj3JX15CV
2V9Ux55u7UY5WBjQIJjcOytkSb90fVss/vMcUfyydvkzvpTIpRc1A6oKw3L64nbrM+UspT5/7vqS
Czc6H6/HQa6z0cH7XMWvsb7dzF+ERJ8+8Z7J5ewqNXT5JKAtxWbn3juPTVns9pNsiKSP63+cn8Xn
KTrS0QV9/9F3JD1AziPdfHfFbPRXCWAXju+8TxE10LNff6m+qfb/M7PR+OLNlHPd16PKkqeiyg70
GkjK/KoXS1U4qLJrClgFUuDo5NZCiZT5SaCVurz4QfhVY/4B1/HmSZSmmDqLlUY6v3U0J/hbPaqe
4xsYnoe8g56CD8zl/dWAUanoRjki1Hu8fDdm4NQqUSqXNF4iMHO4L5qEU/6ghyBxXRhpb8B4sLIE
dK0Hgr+wkDuocUHohskdY2sc5JBgatkqPatzvcSF6/90EZ9VRxrFjlJneomnSSri98ZRZHGd6sd7
CR5PIIyxemLH0CHR0usQHFfiEfJCQh2M3tQikVNd7KLRpcdYwUWNfZ/9iiCt5VjFaj1p0GP13P6m
DfTjgZHr1LElFWY4iFw5OunyM93uxB+AESh1/VGt0sSsn98m/vaT5eLTI8m9TmLIoD0luZ5Q02oZ
oTeO2u6nxMc30Z6jkZkElCh8Of+Su/GDeQ7j2e0njrKh7dpCAy1R3p4pj/Hu0eD0XR0KQu9hpwbA
BWh5st9TABXVJBE6GPqZEdu2qoyp+DHFRY873Bouh6vLo9zvnzlAYQvKGmJcNZCSqDj6YMFcAQLY
BLPKwZ/1U+R1pIeNc4Tjeo5B6IGgOZsWjkUheK1PogYmLlYq+KhqTBSVFgN8ElinJ7mxF85rubtx
t/ZA/Azjl05fzGFcYMh7G9XRMJF3MTD9GPCz3qeCw4iBz9A3btY2idwXClTHcYiDX9BgRrQwQdX/
62HaXIxqZJEbtoZ2mfTyrKQukRyjUta+Rdf4rPiUNwRv60QiVpbkbPcMyzbT3hNMbzdUwADL+K4F
JgBOJ1C1JCaFl7iNQT4f9PMY4tsrQ5gBsUkWwitJ9pS5dgcT1aHePxWv/b9Zv5XeC6pqnP3ZKZ8T
YH/U6s/xCcA7WCy1IiR6oP7gUon8VrSGzYbmTyb0xeBziIrqKHrB53t9vGxp88Be1gN3Npfe0fBl
YwPQuxLHTV1QQcU71wrMs/Xck/Za4RQ4eo5HMW7oSs7ag45bCNrEQV/NzkCbgWI6GpoVFPksrn9h
oKzzaPuvRb8u+yuO9Fe2cVvTWop0AmqTepjTKRXaVmsYzvUsUTQO1rNv4cvOJeCPSjyQpi8+vIa/
cwk3ch+5ZQKVtJzaKlDRR0dZYrPgGi2UAAaAYwFpZBvtLg+HULtvoqw311MRiJe+YZD5VWEtB15x
OZtN1aLzwz36v5EGMw7gp0BZUDoMZH6bPDZmPeaebw2uL94pdTix0Xwtqf+S9a1lekzQQeSzl27P
wLiKKgWUMDtjnhwT4uLpVJmcEpaCr7eCzrOBEVanqJYyhhSqxDKh1PAsKLS/yGhE7wh72W69+jao
JKWMfoVJ2RtMq/4lE+KSr+JceRpKwFTfmM6HHWwbohcKQhRCESPNWCOD5BBJTRkIN0/Gxo3c3DMO
1mTncK07WmuQseQybyyETSiXkGkeD/pJkW59CEc3N2t8KIBzpcijbRtJgevUedaXgMksWqCwTeTn
Q5nwVmlMVqq31Rt0e5xR3ufnB+7A7lwAVgl6COBuF8L65qGs851jV46TptDxu0VuWQmVt6MDfh/t
uU0Hnl0qUVODreMV1/U7zOaRC1p6hDl3UmrA1g5g+jx5ZjmTJYokLa2doop7uVsfjs8ayOzzU9s+
YN7Hrj+daXH4j9kQO1e7XKTFhl0cvzKNHgnUoGNF1zGrkJn8YBNb4612DVwUtYVncOYKAGZWqx29
YEoG0IvhU0um3O06HxK+/p/nyMd1LZidJRIf3GtgXGtrpPe0TzcymV2euCSiDVoCpVTOxBmRrDVe
X7ExIMHdR1N8EF+E1jy6iYPgd5AIkJulTjl8lDQP6f4SxHZbWEg5g7x/ajnOIBdC7vGbP0L/MDBF
jOHNRiw2NN3xWL4TQdluDqPZQXB0ql28fHH1H+PEPrJYiqsVzkJEWvYPE9UUhEl87V5v/BmHE3rL
xnjqvLwNL7fege2LXEMwbkAWRi+6Edy0Oh+3qbxQNJ876ofuNe7rRpMa/PkYEftztQJiWC1skkh+
D2F07yDKFUNIBWdFXhnh224ErP4j9NsNNYUVPj7Wr7g+NxwcEMlUYnlDidnGxR87ldEY9w/EKF/S
mKrKNzTTHjn1oCBXrpmGLVLM/Rx2HOShXFcYgnvxyYSFOpJ3Ij5IEKgYhebnpn/wyVOc7wWZa+Yn
m56n/cgKVGi43W14h99HoeADGl7M2wT8/5KKXnfKj9GM95sxmJpD3D5YNsBVJ3fCrYQcDY2y6GVH
mjYgYypsAtXL1N9QXVyxcyFyoea/bxswNt+AknkfBivj/YC4+M4Q6B3Eu4Is6LS+8FYiBnWXjfgz
IrVKJtyHRv/s7XQSTjy/0ZAusyp6zUGBPS+HlI+2hIvGlb2Iu5MywNrT545LQiAgCrfp2NCAO3Xc
AW/VUcYxavDvusPovsPOjd6dddOhNl30HxlZ+dJZLPlPC5fHnRz+QOrlTfTnL1lKMmyIEoWEgVoP
eVjLR718PMQYkZeXLrBEg3z8Pi4RqIlzTa+DwgeQkpL3H2vPJxUs3MH8Oh691XGmOWmLSqeykLew
4MQm8PjfhyRs6tk6I9gUEHIbuWW7hlwcCzb5BEvHARbIgCINF50caUWPOMAnlkMVqt7z5UIo+0kf
oGNRN8n+uIDMgJKkifCwNvlP209tcs9VZgngLiQB4t/YxHhsQ+VlR6btJR7q0i9ADzT1drq68awO
O+ZtlzSkmi80VEcCnt35nBjJKi1+5AM5EY9112uxvWcDa3TUHarq0KpKKnefM+D46kpYezZJE8IH
/HyEPSvlzuLInSg8gmkawDallaOzUsZrQOJ7o6SKKcMxhV3k65T0BlyC5wyT6f0RD0icUrAn8yp1
ukcF0n/nJnfnH3fAT0bIBdlnF3CqEV8uOVGsCm7+T9buTVCKztp1BClNqJwPyeVqFZ1p/DgtG7eg
d8j0yS/4wxUBW3EnuKueH8BM6kiPIlPFykgl6+Xwj3ns1QxhZfPGv+GhT8RGuS6IOPhlrj9lrG2v
qfR2oOnX8YyQEjIHKaRgob7JnXk8pAIcsAMRCvEszOzpocipQFWjLX+PaCWEzjp3PJAs1+FO0xgn
XPneWRddHruoLm4IOV0CAwUHzxiEepPJ8m9wpJo5vXGfB5MefFeMUe1sVl6JZariH79MrhNBVFB7
EIaESfeDiDvyj4m+Mf/oeQa2EyXGpRVWoXICYaAP39mbgd56vIyGcoYhamhtEnD0MQn/enxU6jPE
VWLpkp94YvexcB2aHK4pOLLkiubDDwxo/6IbV1dn7JtRXezZy88W1j9WlPnl7Fg2R3iEMDLqK4J3
+78L0/7V5bxJ60BwxUmqCXBLtRLtzVDi8bDDEijNq4BiDW9iM/m9H9URcDKCno7kGjeV1EopJigD
7/CZwMRNrbp9CCRcaLor43SEjPhL93BTsOpc0jBIQSEhrpMed7c9geiRhY940m9BRL1omeSyjY7r
6YyW+ItnrW5X6lXEGts/GFITYCdlHozTFeAzU+zT5PWpLRN3pFX3W8ecTZmkHuQM8EvNFh/3kZOK
6BpqoAgKE9sIm1r8U7JFBam0zWYMaO68ihGTmiuz7ao8hJzqq22ecC2HS9Oc0iooXStFNhbhwzvF
xR1S1xNV8JrRz3z5OH+bPrc4jkUi3lAMfd6u1nqi9ERYcrNtrzsklSep3aaDSwflo1PKw0niP4DO
EzK7B1Ile7kAVngUrxw3gIBptJaPHRCc8ZuFdvq3Fq5798wWs7XSSV6TSfkC31zBBQ96XNcOJ1cA
D4kWGWTSGNe1cGl+GuPTDztI8PP3qDXEgclm751xCn4UIE9fIZPKj9dFODkYDrqXrK0McybiBnQF
kuCgDUW4SRrLOcKKy3q09xGMi9aKeVu6NRnj1EgCm92ummqL0dNzHb2+lGCNSJT9bNUmymH+UoIf
snWVVcAE354SMJElD4lZKLClauLoP4KelXgAV2+qskMtqQoyiDdGlLLx9aZNWDlshrhfSLDTEjON
DhEWClk326+FNE4ybphePCii7kY+dfB79E2W1+6g0jQvt24bzchS1XFrddz6W30g7MfQhTsl/utB
Po+2i1pRQQJrOEILeEOb1i4RutuBOv0SgGaNHsitadCfJ145Si5GNJ9Q8cbEL2kfcBsCKV1/DOm0
dYHNZFWQGT/UgoqEH1bxyCw3N6rsbuLPetOm5SCEg+J2RuSma4H4/o8Kl7PwEO3kNc+phIlfmWhC
0XaUkVl28RHc50h9o+9ZRKHJKdWt41oGGOtqIifN2QeJJFBDyu3VCWAdveyPBMa5CXcrumlc4ARZ
heCAkstMmD0itCADi6cVGStBccbwPcKHtxx7kRXo1a+mKEHrB+0Sa6GnvwxtoYbbxEzLgEp7P9kE
pVw/gHYCliJKhQ4Rgwdd5ECMQeXRQ4udHFYwGDDcfqw5veqvLcnNRa1h4ivvZb42g1RdDo2NeZ78
3ECx1iKLjgggWHlj3cfbzWtQMSQIIu9JBHL7nOW1t5Cc2G3mljdttEe5uxGraDJOza7fnPz2UdfC
epEl/QmszmIp/cCJ0vgOV4h/Yf2ND/YMqKi+V9owk3xzvycUfE11D50MPctUTUn0gS7nnBCYMRNV
2zYLk3mbCVe6Bf+jqsqqyNZ3pOuQsYBdFi1Ykdh0CgCA7jrIF80GygXXcS8Hzb5T4gEg+PWsbFsa
xb+U1sBxkUM6aLCDyhFYdhwK11keVBomNbzRuHul87jTK9rS2j2wcMPQnhESjY9GLTIpHTCdCqMF
PCainJQNoJ6T0JfB4tY8wNwkzk91Hs7GWt+9rFHo1TF1zPXzT5orDvzsA0azzFKCq1AD7hcMd1Vr
eMd/V4pvDOQvPAyDF1eUR1MzdD/G/W4eEMf58l2C5LHD/8uiygwdvSGL6/QgzbE4zQbbTkI4TpZt
o+/DxhqrjOVAcds8kXl65FCMfbPTuhM8p/CFFRsvQzVIr1STgUIRlz/UzWbWZsM5NTKdGmMu4/NB
GyoD19MrEPHO2z9nEasKqph/4Go9q9mFO0NvcHn8UFWXPZOGLRMKmDNAntxx/EnP39WFuFGLqMy4
J7qYTpDS0sO69I2ZRGY3NbxPOZk91ayUuX+HlF6Qc5wD2K5/ZIW35dCw89zmYk7nxRSgTBFNHD9E
9xtl1hjNJIprJMyty9MneLl4a5EG6GL5hdQcAfViZWhKX9Ltv4qwXo5tH0SaIR46d7Fe9BH/lByF
9gU25gXgJfGLsfgd3wk4kCS6SRksGVmPz+aGXS/5pXVO4OpFzL5xfFQ6C3x+XuFNtXC2dySq5zhT
3PM8LO9VF40QW8NSOdgNFMiHJeZYnoqbnI+sTSj27EeOYXv1eCQ4E3gT7a2l08KmI4epgx0I98En
7B0QaW4Pb6oZDb69IyfZJV6ufuNOcdEMp2E1V6+xBd/AGWtG7uBQRYcU2ntGSjeu0x1aWGTB5lSL
s59TfdFu78p6rJvmgI1E0iHzz5kOOIi/oKfOdg/8uc4nh0vaikwVbt25TAKk7rxEiI5b/nbLorWP
BYpGbVvmi4ZpRKM3pATH7hQuBdibFiFb03nU/UNF4DzrOqUvjResa4JdBLGJsNLBMuOz9XHdKtdb
Vyky9t0NK0SZ6PKpkc6CpFfQy8W20GyWzMQYcym0wqH+pd3ifdQNtX0wgEIjX/6mwr2wezAlHzpS
WiirzP9lDPirvrWzbNCOKWtm5Y9OzkpfPXkAGape88JMplKcSC+maGFMKKkMDLLgNCnRG8fdF0Oc
koIVlM4YljvrbiTGUSMlXyNBZ2jKGktv//2NJ04eWuv+2pvQaQGY16CzBULpDC4XUtDssb47V0kq
rd+xs/vMD+h6IwtZLXH8SzQz/kCnisF6xXYMpEeeXccXpvTAlrI4FFkaKjFvJfgxw0AqNvsdU42I
kDFk1oqiVvLvtZZQ12FatEGwoAfTu1R2w0kJMjMLKSjcZkvYN/gYMmGWFD+2LMMeQnqmIQZ544zq
mTi+pz7/utdXyNQ0g45zpavaE2vpDYSwgzN3vSiLLAZCffCDKvjF9OE/jNQxBWFwy1GCHhYPnDUv
u2eaR9iNu7K3uLZOXAsjQK0669RAfH1R2eaeEEPW4F+03VosMqZK2zB6atQfHHAnP7hqblOwyQC7
6AjfxPSmJdeIhPbqUGY60HAAnAjVAp5tT/kw0xXsgHfQnOWU5f51FWBezRpK9UMXoaKluO68FzT5
HRS8wosk19us1E3duQ/ctnDbsNv8vX5+jIkoeHXEFWoYD/bjzeSVQ7XpOah1V+qapTsG/qIv63Oj
ods+uklEUNMTpUGMeJIHGqiG4rGRKsIJY1l0Ueu5vkIeTaugoFXK1CC1Xb/MNOO/oHmo3fh8DI3j
CCFRhUxsQzZBzOqUZMzKUKS9dznBer5A2YETREORtOefOUQWzkitIwqT+Fa+X5mxUXLzMPDDvOxT
sylNT0KFXd7c+KxRtm9Q9AODl8Bd6q3LXJRihIZ1rAkUpZeCzFpSu7EyA6FZKc7Ymz07xUvAYc04
zXy5hbJBMI597+fyNpII7XnfXytyZGKVyhm81L+M3XSu8yRRB8wc/eMSj10aZW5VoZl6y5CcBB/F
6cqXVJGoDmbLs+aa7VeKctysGrY9vFHn/QkXu+OEk5VYAbWG+fH8RYSyQgD/N8ILqa7ItKlb27oo
JHu1zrJBV3tySRUa0rOq5N3LRrA9lQMal8Q15dM84jNNVKWoEbLyr728EJVp19bOVo3OzYb9wmfS
WFGzfIaD6T0ED6Y7OMK6pihq2O6I11u8rrTLxcIT3CFBQugEoEM3LkQoft0MusDgBePU0GtlzkHb
9Gz5c2W5rG+wn95bdE6C6gKwfKAHZl/A5WpKxK3V9n2xZRdwwzR6idVqmxWtyRsy9uLFuxNFWCf+
iYfgZMd9tg2pKsuKXyXenIZYQVXpN1ocM6l9S/rPgaWsguQKmOB7vO8oR/AWaiUd8BWJdNN7Wams
VGWoTN8EKGKyUVoFP6PeJQze2GAfNEYv9wjr+hKBiWpb+blfUxMxeP2cnG3owcsJXeafz7BW/ABB
qqru3oRwUavlxsOFjjWTkuJLZYPyWvf2EOozyajkljUXM4CskoXKL8wsFHtAFuA1FIO8mXwLmAwx
77AbnL/Rq74kIPy3f8Fnx6y1AfNzvDYbHdaDo6rnGE7RxOdUmWnMTpqGBLxTcN4H+bojlQfwGdBb
igZHTPV9kSktUCBC4QYYpAaEjVgo4vKWgDrI3JpjUnYPjQoAhwyB19P2d4MPP+UJiNw4hKNOIuiw
WT4LLwdFWLYMwCLB4hl5xxo8V7lowQDfgFYY58MTbDCuljG+teKP286aFtokxHAB+xnQ8P6saQQ4
rtF+tDZ1TF9JUPa3bGuwgSBlzZN8CLouTy69M8y1CW+/jU2/hNTKAatyQJZHrfS7CIMvllo96Pce
pIHRx4d6PBn8wBUYl0+tIy4gHzGu2FKVEXlPQNhtBeyKS7nlXGrZMZ/X30wl2v/PYci/k6RIxKPq
5+ofnNQ90ItKTcrt7LSs4cP6aY8qc5qRBJeD6GqNwOaIRIfCrh7CP2hvCfGG5pEaRVggvd9Cj8xK
Az0+1F9BUyat+h+ei660McrYfbYDyQzOc7Sh4ojSS5egRG7h4EV2Li6yAD0SpdLVX3T+m6opuxzE
nRkZx7eXPrPfHi3A52v4nYMZVUg1/+/bIVFGmKFMfPrWTEXZdP3dqnr7b0ILfFGjIMrRcLCapizO
chpczzRz5x/6CmKYMUC0tTe2AfZP5Iz/L9yPTv3SDdWDN+RNCAJQcD7PXoQsA3sUDwIwvxvq81gd
SI9lqxGd51S9SnsEtUud6KDJXkfhywvTcWUi1qfNDYxNjRrklWboET+0l2QZ3kTmmSpeYvNGDOKf
j0DkEXFoMsyXnRAlPyYwn3UwMGIrutljoQLQzasJklDUwdLT1To+t6mfK1HM4Y7cOUrqGp2C+5AV
rrgbxl8fKJ/O/oO+DoqpaSph6on5MJ0yyXxMHJ8kRwJDEh6va+a/rATsSCpDMUuKsD9CxBluyFxy
r6wM2KeWVUuy5yMd0uyUGIHbtJbfbar7Nb39rKYuc+worDVAcFawXkXWQSlSaNoXUUi2r4pmJE6/
kJu4jwVLjA2U6aX5cXujTfeECzcf3sEERsMxOrHRmRIaeVurb4wlK32z/9E+RKJI0xSrg95hwlIc
gh2MrzW+Z5lPcYdIzIvDaqC0tb4oOVsqY/vWQ8D7uxVagn1cz0SzBFTQuxH/PMV9ggr9kLlPfa8B
VZN4QUOi7AjyHBpV+iYtmBo56yP5Dga3ygTcXa2Ib6tujZl8LxVEItg5+OY260h+5BjTi+aCDPD3
Syw9CY/9B5wrEyKyy2Wcbz+S4KhmVTUPYR7NtyxYI7RcHeUYuH/oGW+dyOzLHaChvKHG0btsDiec
grMIIUsfY753YLD/zCQly9EDHBClvrkwBkfgaHPZxckWgopk1EBY5HDRimMnbWmhqra2bpUT8u/r
KQ+rQ9+IIGmYiHr5XC+HMU2uVER/RWQuZodYcLvwhiC94vDWATGlgNUJLxeM8qKvT1lCThLKfF8U
JPqJnuhC7M9NwC3CVelFwK3GQLXN3WMIUQGWvEYdrW0VejSHHrg4RpI25Ag/7rRRKJC+TZmKvrhn
4YjNfnol1pCiEz9y12fYthFRAjn9cQtPWYUadS+OZoKnp7ZGtpWpl0E0lytUwuaffdefcmqhY9Th
kbe+qAmHyEhhTRv0typaNDTGnmQGOqqjxnmLta0v8qgKrpIXUBXaorm+6HKfcb/DN9/DgXCUbVos
dPrbtGSgU/ti+m+qn1ulLWtWpgESNjl1yBiU1aTDBy7NP1iEeb83oWyXWx8JyfsNYoFAoeFMcPDA
k2YiE6Ytj6wdJx2XlPncvq/aqqyK4r0LrDy9n7CB7Y3SMINUlY5p/1eBe0qeBLHqQ3tY3nTQ72Ln
wj3dfzw43UuCvVe4CWeqyHaiikOXIWO3rjfHI6lHLcA1NVTJLseIsAuvOjWMn5hNNSHTKSjZyyXx
fCuVE6R1Pxt++5fN78goVZ0qlHsphhWMgFhVhOaBYRKBXdzdhrXxfjZ/mjh3EwF9lQZWumRm12Fn
qeMffYK0EXhpD6RR/fXKJ4k3sbgYN6jSlIP0fYfCI6L8ADEoTNB8lLyamscIgb4xAMB+ioSMGQyz
w4WtgAmQBoDGkSqk+22x5sUw7QctX3ClmvzAlJ6n7ohibtfdguE5Iem4pSpA0S6qB7EQrKmenhAX
YRNY0IUHX7vTMqNpbdHDpO1t1tLS7EJlFLrwusgPb1G8hGrhYBcOSe7qnUGmO541roow9uZxaW0F
JEk9EboTC/nucETM2BzdfUUl6SVkcSzbjwkL/6RvXLSQLbYG57rkskQjbETDdK6PNN9wTz/Vl+Xr
fqHkPQc550XEXq4R/Ic1awRKfjtgiktsBRl0Yc7IM6Wg95ClrjdziW7EYt0n0NSBxCLxVtUHRew/
J/CmkYWrKnO4oH6+saJIophCKrZBmN/St/mYLiL7RMi1FtDdEQIlOsusl4WDmQp+jHDdzRTF0NUu
AW5X3K0tzQuJHD5LgyZ23pralhL6jEJsv82TVlJdIA0pCPXEnjJcvH+MgZaxWW0gBwSIupZTPD6V
UKgUkwKJ9DI8rwzSBPFM86KsRrFrSbapyEGRei+HheKZl3cMs/4s2b1D+RXG09T3cw6VveJ1Dhvq
NRxDda+5W15K+ilIw5P4DPJnf675PVqXo1MAdOqpDdm+QQHQinRjJmVEIsH1Ye3Y3XbRp3xp828s
x698IPCD6eGeO5p0zNqa/teQVwYlTn/5XXYGGswtJlmM1+UcmWW/HACF5lQgEuSrILHnGygT2l9H
mOy6GFZpwF+yMDpWDU8nb2nRckwdMk7uWUyit6c8JdB7rQe4WUc6ctzuACKf6UrsSxCLlaCZbAru
TTFtmiLC9TYYQVXU7ulg6s15792JD5+qq9bWHjVi24+g1DRdBr5gLSDBmELAY0LkCFuWa2HjHhq2
t8mr/NeGExXEAf8jzjqioh6au0QZtybns/jdAblvBhtzQPT8ELE7s1ToEyU7tfIKqWOSMz2NrgKB
6YJXDzcw5w+o0/BXtf9q/9bQ6B6r+86n0VNzCUYI35pfka3m3oiMM/U+EDCYX32iPQQ4h1+FSlFQ
WgMaXAKiMgi7TWun2pfaEVFW9wkDrHmw88RIg67ZCceUAlGYWQ8SbU9VLxX0uscWumvIh/z/+rKz
FrH23dSSszWjyWOqDkP1N8dteB4AU37xSYcwkNID3ASslqdHULDqeDbMxC+7byPK8AhG5J7tLmrz
IBeahav1SNkvLXdK1+NpxaiWLJ6ewGHC4iHlHSzeqoc89OQ+zAv5M0eqjIxz2GxnMKh3nboRi0ah
0QoAAopErbwRzwMzlkOBWJEVeCcdKc8JL78REWwiq4m4bGM/kBdm9RM5LVKhNSBmKEsN8QCpyz6K
8ie3vFfAsj7oiUiu8PXe3gjtuj00WjYA1GOwqKxXsQAb6W+jQpnHvQMd91LsQU6fzz3JFoTrvwfV
WbmOEV4xqgEIXKutd7cW6BjJIHTM7Z3vpEl5zqu4PQiAX3B5uiMdGO/EdR74xxDWpzE/B9hmah1L
8gZC0rN4lGy129aM1WjQH9398OkSv/Yedy1gpEV2fal9ePtvBymRh3hQVO2reyxcLun/hDMpyp3j
TemCOpoaEen9kcJ2VgcJ49EyYl2YQJdMjai+dnYGNUZaiyBbrvMAnYB/NKV5gWoqzwh51J4qmN2a
5jZmHuOmHhvA+G8k9GfIQg1nEPDzBmUwRH6rnBtb9dvve8N6g/+pW5AgV3U3qQF7frJ5Ge2sXzwJ
0Hq2xDA2rbhhzd+QvxGJ2tJykkaGaIS4sKXWacABHwT5IeSyaK6SAz6B9U8BRQI7PMhKgo03KNGJ
ErWz9ELHJ6j2Fi32ltCR0CSCQc6pz53B96keG0baKiaXgxe3a1cKbjn/G0t+d0/q8CrjCuWtIFhV
D2ExKXE8z84XmoTPsNaYwlqtwd0TEPkGWqtgc6phvNSWh36wnyMvKzJzeHOeRsp+Ph7v1AJQ/AMB
SgcqB114jJ/9SDPdXZkcmmUlTzR5c0B0MwanQE3S9hK7HSw/LA9xhLDWsAJH/i3ataj6DM+yGH3+
MtXoi0xPmjEwu5F/dIDSJvZwmchuQbWzttOuduNe+cIONlCEO+czvdxQOr/7eiiTB6rIeHFXbSaA
O2tCQ3C8AD+QGbEA47vM9IRgNjVrtr+UzMeMJOH3w9vVr3Tlfvjghr2sJm5IVF9nWmndZHNgU8zu
duywd13rVIwTQv0QjKP1o+yB6jCRGOm1b08SnU8g54aB+b90GIWYQzN1hWIXQTjkTU+TSS1p/lLW
1+vuJqPKI0xFFb/0N+MPLmm96mkNk8HzQbyMOj+gV2VrhIZV8KV9EEu8OFkwiBXECvCMJ22XpMYx
P3e9lVlmRZPxGGRF2wApabD0eRemndfCMjH4Ki68+2C3Fprr639q3OQRkKiE3nJDJ235BzSQq38k
hC87SqoJIG7o6gvA7vtjFWP7xKQDL08XUNAZQ8VCVoKF7cW8u9spB+ddJnbXFrq3wq2kwSuGiqfN
QD+WoXj27jnUp5Mv+oOGr2bOBiReloZNGIFC2h4jhyvkLIilAf5dBhhzpOMGdgH3jYL2kq8V9NbK
ps1QGoyA5lM2MBebObnHY8Hrmn/UJBfsrWM3dHARghnQ9FHAUcaLfHQUT9Iv8amg2YVt7c6GSRh7
o86jYLpUYpSkjCw2f7RS9NJkPFGahjG63HDnGKpFTOdyJKQvzgRDWWSMb2q7N/vbx6958Yu+274y
0ryy3iZI8efPZjuWtpgTDk1va5WG3oKIqYc9YNRyh2Op8g72gR9plI9SQ317EGmJYDFGPC89usbH
hGrU10hYZS0LCG+h/mwvyG8Ym11Y3zCcr4ZcXjC6+6DtnZmtIPoQcZp3ORHYt7OQatIW2LhUy4qV
wv9Tccy4R03q6cMiGTQItlMlbjwsoq802S793O/7JgEzBOyWo6uZcBLFgIcqtAOKnhVL1L5gOnSQ
CCtsLkVcxtPh2wYtXd03BlMp/tcvP3NYmLZG7XYYBqdOBWq3UH0HkcrYy3d2DmsUC0Vu2JIepiW7
SmjsN4kd66Z0OOshiSXPOWkw1d+UnlDjIPQ0i/ExipN4AvSDoPb+N/6mgzZ4zDY+LsWm1+fTyFJ1
IuzASUBc8iY54xnd67rB+vQMFdWMmelZMxrKIaKsiEVCdpP12OuVJlZ9LTER/UhIFDRgvFGEP3bT
Sfzlh4L7E/HLdOXwkkGqEf74Na4K2EJvDvm5RAjffSq5YhEEOhaH7IYu0MC38qmXymBHKueCyrt2
awsJ76/bcI+tOAbTwQ8N+n5nXEbrKhIZfZt3i8tfzFPS0whPPmBVkRL6SvNe7jzRWilGEdOj/q/C
hJ2h6YcKx/IqDLTN5aj3zF7+BARzUyH0eaVTlGBEYCthNhIra4rQ++CsCzx0DRkg4WhwnqnxAMYO
081416mkKsCUuVusde7OAo5PBs4AxRMIdW6bMFqIeUhQSFhyWnWyicshLq9j/O6s76vSfmwnvaKL
8YIrIqq+S/m9uHjM7IYvsyOwfbvZMmfsYZj4J3s8VrR5XJZrb+PngVk3KL9YzV499OT/99zQEBpm
aVBeCjArPwngajgLCGudyIO+XxwqNa9lzm8J5m9ler6y3UfQyhdUodXdX0NI366/sU/1qi/EE5B/
YWXNB0ANX5MajpKDoKFfrAEKr6a6B6h8s51u1l2ljidXqrj6AQbyua/7ZfZcncV7vMR53CsLaxOv
l1hItxvyKNxsZPJe4QerlTRczdwYnJQ6J3v7limmcMhfUJNbYDFrw3UjCNBQ0UezfpLKr/81IfJq
38f5hD2R1rJq1BR6k31Gh3gnfkvsch417Bo0zb9lpJ84UTXuPETORqXX+2AptxPAUYDphOAm0q66
HWAkcqTO4G1k/FLTIktc+xzliG1sCXkJA/7kqs8KPRdwNn/Q9oPJUpD2DbeCwkNi3J7XmiGAKxg1
DNo5HcjJAjZ7b38hZLcQQWnJJZAVd9sTwnG5+RYfj5XZrSTIYYRzlqPmK6J/Dws2ylf0Z0J9+IZ0
1/mZjaKi6eLJ6G87sMmSeq0dLLYSwe+5fGPuUZZRZaFExdty9qihGPK0u+ZWqmlElM+tH6iTLosr
OENPFSR5bkFFa1VPhgfh6C+3WSeTxMa3M/ZIZ6tDIul2rNNFfFq/k1ZEMn+lkTXHAGT80D7g1+m8
IMYesbQa8iOdgj1maCqctQCcin9uM4MMYUhmWkWaai0PTxWdmPEvXB0IgR/cpesJMiRCvK76ko/r
ESopDaEZsJlOrx/DeyqRg6qenS2eBRpA6MtPIUzF4zSkYByZllUVxRjLc3Zit33g3m7FHRTn/Eeo
Cxn1lTq8i99meFnhkg5or0Kn2mi6fzqR53DKWr4dgruRyJ7cPLuD/IgKzND1kERGUmPZ2J8Pf2h/
8O+J5QEZ1NaaeHFPfBAKaRAcHGdenk8/ZEV99iVKyhLI1lZHcqq7T4MMGUaTjWVfgcnMpHRw0vB2
35428AlrAO5hal78OKardriTyoi0bZ6trlfs8ZxBEjcR8m29p5nokIeRq/m5o7zyfg4FFgXQ877T
CNlFOIQluQ8wridE3u/y2/faGY7MfMNY6gabzghiPLR1bteV8Dus/myLlxose6g+U0tJKSejDGfl
v8IUR+H3erbZQR13/MOmuueOo7wRkGg6XIIRak98VSgYfp2UBTgIIcC1QBhziT0ca0MUT7TlaVNA
M+2CgUl0VsDKmUw6ZlCGp6K7fc9uKlykeRXOK0OUl8vcS3WviKWagHLXkVbcq8edGJqhAvj4GkRr
v3CyT1R5pxwCEj3NGuXy+XX9Ll6Mn7qlzZ3WS2pjUICg2dl9GPRV22USjBu4tNDFsaPXJ10ucHLA
9rKPk3ggMzhp0BFgGKE1UI+GJbJG1tbDvYpv7rtaC4BgUT4fhBzEyAuBzyurlklEpNkYDpnn11yP
YhiW3L67lmmkyWpA4SSL1un23OAYruPbXC6Tb1u18YsZ6rZatDpumCS+32s9Fk4yQXh3t4IZsdUJ
7oe7YguyaDSoy8ZvgjSBEPcvnNciu8Hu4HCH34KSTl8G+3LjIAsjwi+E97A6iL3LNxGaGdfpZsg0
X4ujUG2wNcdP5mk/UcAETjaSVApRFO2+2BBAc1gfaore4z11c/3Iovb2Dhigiz2TGKEcq1QvYBkI
UTdLXjlcO5M+b58YYdyiHoEkpfjleacW4gS1J8avTABDc6zDD6/ZjN1SJvpgyH8GRsuYUELMBR4S
lG4qtCCmqP3kGodinNlLxUN3jLON47S3CEjtoeW9jW2r3TQiMm3o7C+EkWR29wuBH/caqsbDozph
nsZzixPLZNfUlwzYmDF7YqZTcQbiprli0l4OKgLQeQ+/tvkC4hIz7QHABZ6yk1ihr0Iqs5Z0S1K/
oQcD70a9sj1lwgKoYUFeP3lYb/Xed7edZKYiuz7eD2SmvYGiKfl7qGs+jA2RMyjRc/4KgKyRM2Fz
KYHAzQUNnrrFS+PDvc9u8e4jZqL6vTrl2mCkPmx3NBYxCJJrSqckMAVRDo/OeIvDfmb7eilCoscB
6MMrdSbh6orueJquiT4L2TzugEFB22ys8OIWzjV8H8gh4oMgEnJeI/9m52svYAUdY/iDrv8zklzv
1dKQfbhjiD6Lyd+23MLNkEmxyrNrRRN3dG3pQqXh1xtISVzv98KhFt3nJ/Vp3ZaQxs1OH5sN2/b+
y61Sh8d+3aDG0cw0fvBUZCSFO9hGa2WruFWpgvW/TefByH9Xv+prcNnjunPrkAqRSbgCpgE9AoM4
p8gdELI3gJ4zAesWKkS7oBfD5hw4oOAp+u9wWrxaQjPjpqDsOEdQPmQLHe7Q8iRNoGE8OgWaoaE7
FzgvdZnsBh3+fzqdnZXE155AcKWuZ6ysXIkMMyuWvgJqPM7fUN/4sQCamRKHi14Z6jxjh+MBRL9m
xx87iOsx8sTZNMnWPzdaOjMru2XT62HrS9YQRPRHAU3ooJuLfqgbuYNSX95c31+QzRGz/wBCM0xa
DQePDdVC4m5OXUy0tws4RtJ2OQx8VF1g/6p2V9XWdX6yfS4j7Qxk6v8ni/xl4MxY/KJT8hyem7cF
RDO60VHuTNluZisl7gQ/Q4Pf3nF3SNWNgzNVcakPdi2pKQOGpIM4jiEo3KS8SHpOtBrT2TfvBCZX
7O527vXGvzKNf4+DbNDzxtG6JZQzlCF6X3aygL9nLXQIIWhLtApOsISKBKP3oWr0rMZQ0PCuQdFZ
tZFIdHo63piOsZTbUJd+IssjiSqlaQESOcjX8F+zITD+MvqVI8BmZajK9q1aIjhx0XaoXoPE8jOa
6UYThXKCA5+pbZD7lkAPVR/pBLtHrzX4iPHiEuUWufWS8IjP+YNYereHPeINW5X0bwMWfWhQnZAy
DePE43HQBpm0IB/qCvQGl9LKi20/p95Q9w3FwgIPwr0jyhHs8QwIHt93XgOyR2E0K28QYGvQqyiU
zGIVrVviKBjoE/lxD8ipgiFAVStmKV1GsZH/1Lrcb0XK+D9YAn2sDz9EMbaGOndYipqj67zDTQ1i
CvYOzlca+vTFMGvnMn70ZgTDXFL5rsS7bbPWrWGPtH0cmrhhUrl02baq+/njPKfUBmrzE2YsyX7v
ujT7IsiYFdzo+P6rZX//yQq0svLvZfaKIZOjDPqQioFtrxg/qe94uP3cp30Cyw5Yh0knGXrnmRk8
e/22v7bLd/8iD3CiiBHlLybcjtXyNCY7rZk4olALniv3Qrn0tzw87TtvqBlMDY6Bya5yrGmQXwI4
Ft8WhUsyL/Y81uFKhiydvEkWPSFvLdiUhr+yl295MscMtfuy149gsbDJIXb11JhSWZq2XGyTeMXM
UNnEAnz/0HwaS8kT3gmIR+JHuJQg73794LuMA4sxh43FJ4luDtkSZ9PT2UoPyM+Ih4hxe7POapEA
9YRsrlOOOPKTMHnt95pvdWFTaHZndv+rEJ5YnygI+ERyG1N85SAaoWMNFUyMPdsJtpProAIaObMg
JkiHVycudWuLRyQq2LMBxDi2ExhP5/7+3o8nmQI1etqvux6ScHzJp26+IUDlyv9H89+LLSdTzTRs
4Pkwi2qsbn4NpskOgsnyUh915EmrTlzw8iwp6GfpAXRXoLe4LVJjutbbfPbdLMF65sSLpRoEHQoU
NwHwq/lr8xSO4dAPFtyto3Mxmq3UzFobP49PEn0NKi4ZmQeqcc4W/DbxLPvJaT2M723nLW2zKf+i
f9NXzA9QJ/ATND7MBCZXD4/E8DvNVLdJgN2BrQbB7pzrmQBzMBznOoSqmwSIiQRTzKTIpW8EnbOi
LKcwq4u9ERl+roKUTWAFvbnWt6oOVuQmRLFC+7D9yikxLY/4xlhzm9miTJHebouAz8Cjztdgaior
cUE+Hfi7w5jLCEvfHS152gLsO6Dl9BSxPnRWtjI6yE/aB3407JZV+nPn0HtsRmeQu9rYUkN0sDyf
3ytd36KIJ4kdnhPTEkc2X0fspx6SqO77uCXr77rbRimFwtHPAKI4P8IalCfw/RIUMJeeuAEs+dku
p5UBtsnPUnwkCF4BThTdfAV9oz6255UHI3QvLanRN+7MnVfWLevnlPgT33wxpPgJvlz8q65WGVxk
5cfeHpMk+jx0qOUM9en9RkFxeVM7Xvo5oaD3lLz+xXNQDhCskLSAKVtsOuf1ngXvtrL2OkAGVaok
bp9GCSAaOos8TxCUM+1ehzGPTjGFgKDKUsfP4uf+GTOn/jWqmW4Z2rqxOM+m0ODuqSh1IW/ZHidG
HksdrAlwPILMwb/8JqOY+W9sXO2xnX+/9BnzzwxUoSuz+3ydHkENIyu1vFRZs0jXUh0JS+ApX8fa
/HM3EpIIcDlBOAXifOAVN1Olbysh30zI/5Y24b3i6DlKzSsBMyOEcVgbeRH6SXhp3MeHOd4hEmX8
eQScCyKDs1QVLf1gSq7QdLkgXqBgiTrI3XOfqnsfPi33786xc0pv2ssMqFWkBgysL3jf8hOo8V1J
iPczVyc6eXVercjn8eru8L3tzhaEfDJ7QDOoySAPhn/skH9zTRQQzidItkrub1N629CuNiGPF9qf
ybgjcJsMNMBewaLT+qaWfjLUsQbEC5sisRCprMzefsDHs7Ef5UgwOcdvaheV0zSCDjSzSJWzSs7r
tYhZtsEldvwnueUoPRyX0vg1C1BaU9KjL1lsGcgAsbQF6rnutgEsgS/6it1cxiGhPCUDHQw6xSEq
pE0valgo6x4XYHNNAF7/kqxU7AY4fci2dYSW4+jZjcSyJBThVbTNG3VsQOysSJyRu5yvtzEdz0QD
4AVjP3eyVqrsaQ+PZ0bjYJM1dg5wuwKFcg5gA1eTMF7nCwdsN+tchFI8X2GcChZXEknlHGn8JKQy
1/EMOU8t8urJIBdM3Le0hKyNej0ORWYt5SHUxUqXLxaXQLF6/CjHzttq4JL5b+AoSdxKgGvmbYuA
sCe/qOP1/v+zeXKReXtAH2tjGr3N/eSOt/LdGtjWko/Y3w4yRnqb8O8CZYTnrGVMGuWhjefIOkkZ
5msE98CKy2RTLQWrEcDAaEU4Fvn55yXpFChyerSxfKULq8G44Rkg52vj0XWoOlK9t8Gep3p6YzxN
r0CswOBAbYooNDwkVbjG0I5o6OQ7tLqTiMWLbKeleVJKizntrrqD5vOvKKU65X5qWY3X2gxVUjty
7b2l3LFmwoxeDpwf38rXdfA45ziJAiZMOk+1cvJi5ile/ehfMUCVzAD2N/cvpMksl8Cp6N57xPWR
RW8Jyr/VEm8xufJ6BLyFo5zWygCk3xFfRsLMvcZUBRy0cYs7ZaLLwcaY+koxnu/XiChEbVDDDCGk
tGmrUBKmbXiiYoXb6oxDlfxB9Vr/8gwtausrWEKBiK1Uuxaf61Yzez6c/rlfBocARhFU5WskhUkC
SOwHkqUZyu3twoEH7Od/GXqkakVTIH/bsG6+NVrbp/Pj1i44vvmyF3A1vG33qLlD4gFe+wL7GV+2
USAVQFz0mL8+A8u+9XGr5rKz7iHsCAoJeaTPYSpspK99/IT0+XXIISWsU+U1NR9tp9jBcm7ulJUe
dSpov0Jot/d7t7HJ6EwdSASfRmg7snUYqejWGMGIV0E5LNcj7KUxP4qpFOe6ZrHtrwhNgeK+lSOF
pdQwXsFcway1zlItvRT6Br0tnVnRLSt60GxccMrn0y+yYe04ufe8Sk0vSBikkAQKg/gnrmLgR1yi
VO4kwXs1rWw4otn4rExFC7lTV6q1xGaHNX2rz89BwNdYMXyZz4ocZ0AxyiIVDb+o2peLbNgz7l58
tHrhMB8nqJU1I9o4TsPskc+045GVFEakiPVM+9kAuK80JSFXERXc4uJdIZqvJip3picoxpEYONmx
1p/eonS56EKwpZytkH6tgalPYJyjvYDz5+b68QOrfR5licCKazC/GtcwncGYKG4UohaH9X/f/c3t
UefsStNAFKDio0+2/hcZy3obgGvrEAUDnygNQO+hsuxrqUNJDTt5fWF5vBrlgHAhqB2vww8jZMDv
/Ir/wkjymezWo2+4rgFkPY2aj4ANQroj59AcIzRkXRZun7Io9o8CWyCO5Aqx6PJHqkbwsZebCCpj
kWhCi13AeK+InFp0XF9Ic8P3MS5lKrW/6amr5S7FrStuOmSzdrM0FFXEPSWhOY0KOPHmWIOLIoMF
jGj9DmtIChJJsAqiulYuq5x0VHab1DB143vw0W0obdKqY8i7RO/mi22mPJ0MALM5JWPLLTqu32p+
HHNeMsEgypdSrzv6r12DYH+NlksRz6mN2CVvnv89y2THPRN5kqCC+ZKNaXcd8IitF9jwSeaua1Nv
SF/jmo5Xy1t2ciG1gL9k6ne2PeDWya9avNXss0Azbi+gEUVEELP/dbhQ3xdxIgBA2HzLFmt53fEN
W0uVqBMpJa/P/gmax03LlAlVIzm/pvPbcXepuz0BJ1v7UK8EGioC33dFflyHyv2SzWh+7FU9Uz8i
6gp8vIfov4U1iKQx9p7ZNDN/bZriqf0Jo8i0Tpl9umGNvJTZokljrLgdaqyw5yRVCiz1Way7KDiL
JZP1OlGiAvunintwC9fQLknbloJS2ztJNo75pBmQBGPha6UxowVgMW/NiAZqkdZl3M0G2ZGpobuc
KKcZIdvq3o8zsNYGSwEQW7wrTaDb4LM2orLVptz884fI0p198JbHW0jzwCc+u0JjdZlpdpQa1USU
6B71JCGqtHV9t6hMEVj53GgFYhYCLBqc8HBwkIOVeyUsPkAu2jqBGs4lY4BoHLenXFM4+Sf7EOrX
s8dNMrGD7srsnKBMP6yOcXA7ov4H6T3bF+DR/AIAbXeWd5IKthNZC0YxGS7YHVr4gUtc5Y31RJeL
XNAg5z7OYZ554LtNzRxfie0ruGX+wPX22FaapEJYWF9GFzMvNKIWhkKdGvI6tSjDSzl/mbnm2jX7
508W2TBmG2drU0LDKXsWTNea07tbmJBR5XAC27WZ4zONderbwsssBBpKibK02V2MCRIzttvgRdBl
yYa63P3CAqIR49wPChrj9eTb4Y1n6ZqwMJfeifQHI+lgRQnr8vz3fmv69myz/S5C4dd70q+n8i8S
3g26sTtghnvip5joX6NZxMCNpX8ngCTS/3Gcnqm3W4FKQP+F0helAdoEdMlCa4Fn3ulLaGI50x4C
gkB/jrUwea9hqU/WpIKHRkXQXj1MMRhw6ypprIu343ivnPax8JiNSSn72N5me+deP9akPeHuQ2O2
wQtXXeBGhOyPSmmcZXVRHHlv5GwX1steYsNeQP3pUndvbiD+18FG3JX2bmJJgETYCqmcATvAoPsz
WqT7B1e++qOwFJ5JEXGKC1G1bOlt6RRoSwvo3SiEgfYLyyBALIhmXimV1uOVRK27p0VX79dw+WV6
YM3q1GAZjw7Z5mdl8XynWLERPfY78R0BYINIYlhuMGJ82t+GZYOaO0qvnTW8x+pQqzRrdltSBAy5
5F25TL6m8ZigB1V+QDmXfORxgQ1ITYFUs0esT9gmSV/D23rVIsJ6SwLUn7XQ0Bq7gdz/qNzxekqS
raWE1x9HuRxNT+yAhBvTpc5ShSRz9/7QaWWD3gHl0ih7CIW17p7dZgFCBQStu4iV4CYcNRcHO8BS
UH0ahFlpVKgbph9uret0ifCrrT0fyc3EImoSv9zmhDtevj2hOLKXf4HO3i++p5gqARh8swcH8BkH
52q3ijWXkQ1Vly68rwLbksbci3KJ/O+2UCz3fYdm40VdSbFkzf9PB3BUbAQu4um8bx0/Ey3EBp7w
yAwTF0qMndcHbQElawW1pyW1JkMvgRfBQIzn4TcBsmmNbKbQScgRvXQxitthDa0JsePnluLQk0iw
qC/gsglwiItWsMUjt3nX+oGqN9DXvBayOopY25cWOZYDvnauQ+DY0cb0ngrWvRQyLXD11acKS9pr
uwC1/hSGncQFAo5jFdw3broHvrX2qBHikz3Fo3vl2cX1ihz6oZl151DYaGcbmqBV8wFaXGY1nLgp
lNDpoQ/ds4TDuIm7fJWnIwuP6HptXCYuqssIqWNILMhrBJj88zB8JzUol/4QEQFENs5rLZnb/hDt
VEVrCA3ynWte/IjxfGIaQQHpEH8nNZuoyHx6ZZ5AJhezFY+rXo32eg8DXlFVwKPd6necb1GXEi7T
l/pBBokT/DUQaHAPbtGl5Hi3CEy+xa8ClcDiS7dR8Z85etSIBhsJLVHyuX6SEA7u0hq75K4EQFjL
Rka0vC8dHw7VI93LliOYo3rpkFm5aMSNevNyxYY4E08lUdybiHRZp4f/JOzSNQutmKi1M1R4F2j/
NUlC4N6iH1cjFUgpIGxwjg5mzvHOlElzV+Oj0P4/6Iu24gDizTt5mUqJFPtVopfMacI6K97SicH6
oK3EPqFy8pFUl2KIIaopuYrfz0pZer9RMA1Tf5JCddULM3GvhGayL/yNBnXlnJiHleOintVUf/rR
HxyImzHqALmHGaOLRRlvuFtOQJ0rT2eD/He8Yv6S8Gz0d7+8SIWaDZ0stE+u9BifR8weHSeQXNLw
DkgrpuGq/2u4WdVjj7bUGIGkQtFouXTQenr3zpxteEkBjLinPa/dLBGNI3myszAgA3qlu2ynlc5U
n17MXV+lJG5rxctVY9+/+66lftmBI+xnLOAm03PEeCYfQGVoDRxJfl5TOzCrVqqM+U+SFzpH2Wx2
9cN24fEN8wdWb03iP9IU+KLEzgT3UVIorplyRFD/sA71DpxuteEvkYaypE/xMroC4IMUq9KUNFSv
CLLNcab18fm+SGDebOEcwwiemI9Wgbu53aMxKDTIXPlQUsuPboQvEc+UGstJjLZYSZSXrgcxmrGc
wTxD5nUxWReO33e7tyYc/K/yo+KqdXDJjYrSUcDnlzc8gK2nhO4U0iLB/SMyrV2Omf1TuBcb5GlD
UtDrhLJcRr4h2JtxFDjfJrxHdY3Os8VO5zG6O/375VnwmFcRad8SbemnRnMbCkrBZOFr0lO5Zkcx
g9KcmvWzn5L6XVmXCRGWAEMevlCdtTDVJo3/r8ysUkwttRjp89wu3nHdQ0M9zK6RzKKpvspBBjKn
MtLqKr0trJ3DOiqkptE67wm6yUruMvaqCHf1ZRe/mRDoHaq0oEwpOkmZBqcXfGctIF7OAiSxBW6j
yoSuJi1bUmbdjJHETDYgSKKazCZU+NFt98cHkruIL8J7Tm2c6Q/WqRfajr2x5N1zWEFIAMwCxMNo
UNsg+EumRll67+P4PvFGw4yAbM1+GzFg66NpzB5bZ37JHcxB04WMo26MTjVXewPXDRMekXQ5Pen/
BjyCWbe0NDsrTABCQYy+id2mh9RN5uMcJCOl3eIicQo9wtk/xknmUazswqHQeAMQtcsoYTQxymMb
JVW+asYtFO6h1tEllNv8FS/SZqU2eDhGfrfmd7NvFdDhiTbnADgem99tpfYHBtJE2u3GzSABB5JL
j0dnXvdlfZfW2CbBzfggqwoQch4P7600IZNFfLRgW2eEuI+0SO/IiMC2u753D4IqtVRfnK60nDW+
BKcaFtAIt9ZMNMGPC10xuINs6oogk+9zBTVpPiEjpqT1AUjF4v+rK4outwMoDj9Nh4+qA8pA9u/j
/7tyaICVsvwttpnMysUM7+xbnki6UXv2wxBcYIRdDSO04lLfdGpUrVrHAiWHLb/KDV9BAEOHCIIG
rOUpXLPy9rhty1fta9Y9SYgqiq9dVes1GuSsCBEFT4L3Nkhzuohj16quOwcuZ2u+pBnznra5hmM8
cVN/FMsxhtNGZsuvtZDl1ONYHTDcLo9sqa1GBsrXRUt/mDlLB2CzvxftEgrtxAcqGZ1dgO83yO04
0s1IMZTD0IjXb/qSSU3CjUSRhDXdzM2RYEfr473JWJpyRefxc0KrCooHDGzPe8keyQRXb7+bdJbE
00ea6l08gVVKGeOrHO9mJk16vA+1K9N12LHNqLYHT5vPWF562ap8jRqAbQnzMk2L/7ciWJBP8QYs
VQfA875AHJDFbwC/QZ1+4vjdsqG+y1qIpckLvQ/QNG0Dw/IGEjKcaUuNUhtCehEIF/Eb46hkKR66
Ud/WSDAtE98ZbkwXMJAy/2+IN+FKHPQf0n9xNPTj2tnjmInIZ70xFIfCF5PXiKnctilkxpUpVSvz
GtQ+VI5gLYzneZqiD0gvxtSkzSTMZWF0znI4VM8+9AE77g864fMGY6PBbvDlSCHhU2mbVbZEvL+3
UUhJjwkj8QxkABw2NcBzksm/lCPrcBpb92gnZCQB/ATwy83Jt+ly3gyoHMInQ7WEJS+vURgyyO4B
gLdAx2zPlxDFNGTPhxhE+va0rysQLFD/zOr/HfCqnPl0Ei7dYSRyUahVRYwaWm7kmvKC1gDzTz5q
67EU1ippSFT6g9RcZfU/4Isv/vc6Xpn3pLCTu8i8remOxcmfeijuyk98Tdlc0Lin2m8l5M50wUxN
FEA2SZLD+lyIP/r1UBw0Fpqy50FPgQKPo7jaqLYRYkNemUDSTP6kOH8PVQDU5+gwPL6H/w3JKvKt
T9qMeduk/yZXw3azfQd1WPuPSaQTt5/lHIS7WWioUJWf2FGUQNbkxgXe5dj+85R8iK88CKOb1fb3
jc8h0asPq8rzc5Q11LmRCR9A/Dw/aC9S0ZP++vPJsEe7Kad4ltvX8tY293vl+tUOOaRghroG6hWa
yd19wvNAU2hzmF2ZYqMmeWcwS1NrZ6PvGtkDA5vse4QyiTe3tt/eQAkSL6CLeS//YObqKVeX1Rml
L/jpeDKPY5nPj+bGwIfL+aEOT8MR1y3qIWrw08QEVxTLDbN7/MROAV8f31+yD189IO39h8/wBYbL
y2caczHs4qEpsFYqf50ghsQ65W0SBTCtqTqFsGfZNOVBsdPmpGR/8HM/OdkRwAubwsQjPbQ5yXjb
Q62GDGvC71dDf1iWKRAi9ewO02Aev9ImBIvhZZsx4jG9gsRwtYhxq1TL3dyGddSFzoh6j3rEMRID
w2CLYuakHSbRd3V4VMGhRpO45SGPEM6vECeNVNVLLbMByJ8v8JDs3XVrzR5tiDgEzzo74cdwSyf7
pPnpdVUOFEJa2+tJsBAJeAY40oh0yY/FE6Uyzn+b00SEzJ5hJzvK32nMaxy/AMtmiea2MuleK1K/
Smp7tCyUcQ8E1IsIISmbKIvcz8p8WrsG9OKkCLgEXNZ1h6j/arI5zd7EtwgAscMtwxK0ROL52Pd4
3t5SIoSAjQwLxt/zT0lxq3SyUOgQA/tyMsQU7uuRuOj3CUbg99saPmOug5VRfWcj8UajX+/IgY8s
zOBLF1qa+G+e3RZ+VKZ1ot8pCapd1TO3ESHYwM0cgijUZp+9k+RdtvJUilBetU/4FgfWieKSZfRG
E9XOdaucdRss6q6PzqR2DT3NOI7IYat5pkJU3G8oOoUQ1yFzkMWL362CKiMe3h5lqgERVzm4CeCO
ood+I5Hdzk7nOtStcj7wTTYBV1hzocNZam0s8C3nc2xALYMDva7WAt4QWoPs9BX5i7aa1Id8HRfC
vI2t99EPIvlplmIyef9pvHCOalfXNhP6my8GDi9RNljvzkn8/KUH2Dc/GwwU5onTsQ9PaxpVjIu4
g3k3cRzrbu2eHL/eLL8aMhJxAzuWlCBA9HfpakLPrNmGjjCq+1OAVrQDwEhR1BK0onHaUh3BDg/Q
rQIUlupPnII5dQWgDu3rr53etUfwthtCk1fKECXqYg1+7PUnfiOjgD+Cubi0Wr2pUxdyk5ctof77
qG/62TlWFtYyG+yITSrk2NO/nHnz5HQHGkQX2Tc6u3g0RkVZgbG3+dVu9f1o+3gyoIR95YDffS9s
fYlJCJb+UaOb0NRyIImayHMfRJHj/2I4VCxAlVARb7eZESIGbJGNym6pt9VNLJV+PJyyGxo1Mq3R
TQPsEkIlkQDmEeX/UbPnBkQQuQ4HNMJ3HdvMo4Eb6Cq/aIB2aB9sB5BonSLiH+irJGlQU+jo/Yql
0bQ1VYs9YIaOSGYCIbupEPlhc4r4+MOvdmaGpwQPN//290PWltr5GalvLg//GjHYeTY/lNcJNxJs
K9QoK1tyOpBng/bE0C84Y99SFBVnXGMLBUAz6Qn3WKnvfvRL1Ugo8/30ugXmqw8zv/VRTyRIJCdC
yIXZDjrxIXIltRfXppugZIdYNMxWhLggj0vM2UkS/PkVH9qkJ75T8tpD96L6glDxvJQyCS+8Gcf4
cnduQVPIv/oQENuIoxIbmSJj0LriHffkJ/XXegq9fCeA6E0hl1OljGBip9s1F9yCGtLRsXlf+q4k
lZjuzTRWCMVBfhoK42O7y9S38EpXMZAPCpwa/O0MU4KnhWYVtXr/jlAHJYkYvoZJT4J3hAzZlkxE
tOeCMr/mPY2XKBTfx/fQalcpAj87AnTWkPrX361Z15hC4dZOs63KRuX8auHRg/VStf1PYMLOS/CO
8Lfv+fdoQvc48fxsPO7/ola2xP8XWKuWepFnPs48+Gq2GBD/anP03JagdXNQvJ9nDpPpXG0o3EDj
GRbIJFO97wUNRcGCKF0TLC5PuiQa6z5uLnnvQxowneeLpnDaxCqHTgXSoQzId00Ii0G4NXCVGn9f
eujZjAcuuEmm0GJVGZjEgV1DYbb1ejT4A1aSkhk2wMf+d0eJmsFtADKxNGivEd7+WPmFCwBWpNPD
mmUmE7KFvE6GXLAMd3EybyKPCqYHS5WkUUfTtChvSm4Z8PuVwxW4sw14MVZYUSUzPqRK4VxjJSon
Lo1VvUBETBRK9111gVNKLFw1o8sQQzfyECx1erTpX+/C0K4FeoM8q8Iqkc/vZOkH3wjouRj3ArFS
C3RApKJY31FWKnFEGJxlJ2/QAyghLsAiFKzlwD+eSWYI2vpkC2rlNgv6xYHwgciPTxJWLAskqerU
niYLuSjQ0X1BVRZl6h31Hhr0Q6trJSx81ucJPud+Kd0RyEaa3tHPCvMV/2WnYAI0DJMxrkWzA7zx
fhTRTjohDDPSftUy5K367UqQCOq4F/lhwq7EpAVWmYuYeKPa4DLvX2u9tya+JWTL4Nz8jSfPZJ/3
BkQnpOud9kydEmCqJS8zd3XPo4jer74E1po9ySfCewmJB7RR7uQ8QwkR0e150pg+7BGb4YMifghh
XTH+M3006CZeqrr4zjnGtpdEYFX0m2W9sw6YzXWVNuaVUAIqf8OzBDb7+JOrVBmi98TNmYA5MN6Q
CBXsLL7yhlDSrpYLWegtCi1Xh1jDC3sFlAQG1nQo+SlZpRqrWFpIoKEgCFWflIgnja88NRkQGjWE
URMPQ115xO+BYKkQrxfBmfYwModpRLeoFDVO5q9xDUk5+TCaKH7+kcYynAS1+AiQnd0obfwQYCaV
YvFG266v+FIhRamSn4WhojSWOs1Uff+RgnzzEv26HK1lbFl87jwjf+y7djm2Cu/EfTJlLkSEj4zK
2UTpoNQW7cSrbmSYVwBWPpuwz+3Zdrwhv/IQAS/06UDUN54gk5SLlNQTWAQzb9p8Vqoau6KnbNIi
c0cWxYxPTMQenXdHadJoo/BOSzBnn7RQzHOGQ6adN4lZicd1cSplaVlyIk7JEqDCse7KxLDjO+SC
0YJRrUcAOKSkPhv1B5qC5n2UO5utBO7CwVF++17pAC1bC/gJ3lLOcADQ83MFqMLbT/ovl73tX3Ok
x5BfA96Tz5rB/n7ng0qvzObVSm7xW2v8EWslhNz6rSYU62qBdBjWztrjZ7DxOjZU1+pGe9eE/SFE
5aEW9gg7HifNM1p8U0gc6HiwRJ9xq326yJOx39hcYaasxNExl9G29zDqm8Pq+Bgs/6hNHoWPCUhE
MOBsX5V5J0SpNfrErEgvuWhZq8srKzxFNVZLmFMIoTiIOeXZ1+YMZufDiLBXnZpsdQ8BqUuvFuwq
1zUhSmuG9yijR2x0BhZy5CvsMzH+SUHSwBWPjQRc3ahfeqXorwOsdWDc/4x5unTJkEBGamCu4tBv
2RDBcFLxp6iL61b1+zrA4JPZwfntYgeWJfNUolZiA/ycWfwJgScKw2jYvBgPDEJlSg7H0qRJohbT
6lb4VvWQ3LzxmvKt274PvNjWUPVZ0wjBhTKb6vToOl9a12Wf5yLwHbAE6JfKVSwcc59oAs/hI4r2
aRLDHa5Qsyegwby/VVsWZxR8bqeCuOFuUUyw1SXL7ftxCkiP0hgJi2OnTKGHCBKOpDEcf8UwzhPx
kBLoafdYJxSQJeXOlXetEnf4QFjxnC2ymnPuK2kSGs0Yc+3cf824Tt7QsWJjnKeYIVd4VAZQz8A3
nttL6e3dWAxsJrZjpvUPBTkQt7P8jo9QzZCsla+1TTf2O5Miv0jM/KSXTJ+w/WABwxMepkTm5oMH
7//4iLkQurFFuc6XuQ5wIMhT+jSpZEYewlIuFaJQWtsmNxLg0QdGUtACWcndS1hZp2TuJ7h4Cgqq
q+pRIHFUeVtB8mfUmujcK9Xn8cnMb92SVeCaLVofg89K63Cy5+AxAPuFZwCOTb3lph7fa3kS/St2
YfzydTuF8Etq+Nx/6915dtsP0N7yDLT2/WZ/soZQd1Js4Fi+am/gYZWX7x69gadgpVei8dlm3dAP
SCLT5TGsnUcCKr5ZLNOWVroqaDQKIlJZSRjIne9Hr6fXXSgd4OmeL2Q5RVIztsx2rlRpPZuyf8iQ
xouDh4YfKYKi1htYJ3Ih1G8AbF2pk0B0334p0kvMK6qOo0g6Js5SF1GsqH/+lSByDHWlnza0Mzaw
x9UuAVulzHL0AVPfCygU+JcMQfzqg0W/CcEkkoVFt+uo2HLg+Maw81g8avXYyijcNgbxoaegfvju
Eg2qIxRbjrpY6l0F/NIQmE1usxtcTXp9LkXBpAhnjJ6p7E2ij8cpESCZ05KwoOp2P/hBzVLaqvsX
2BFo6fTTndKJKJKL0ymb8X9RusEPCZgfyJEnwVYDl4jqkURpi6riyIWp+Oi6Tvv02y2Grd1AM6jf
PKcadTxNMdS7IKEJPzFPzsiBXUOk5HBzO4FeQAaR5CX/iP5oBeOxt38cBvCa2ZaxJo5JGWmXsgyL
9Vu4+gg+0uzhnQDVxOYIB7/HljhrNdQXg8UxQ9303PbIOm4gDNvyxW63aWtebbR969Y3CWS+p4kd
fnhvK7RZHgFV/cxH2STds17vM44HMhUUvy/RtsQ0YfV6njeNGptA5GUGlLmjp0UPf4Bd1jiQjO0v
2u2Ndq2NPcrEhIceiddlc3IniYk0J+amTdsRbB/de1bh34rZtKBYJaxEKyKPM+3g2Pxo5VAJkOAA
stfrXCp+i+T+GsZofl6hdCBgGC+XZ+4TlPTGc0Bt/eTKpuHlWyLaif1Doxxh9ghOcGPlOi0Q/YJX
9wuH7ad6DNahky8ETOVI+hd14ENNjTC5b8oGbzR6+KjzyL5HFU9yuGu941GAef9a16ac0bpSZ5Bu
rSznqQ233YJFV7sGGMytprySxNeXjLVCacBZyxl2xH0zeU8pAs/AkiMyg/b/KKlQagWCk6F5GA4V
uU6kgwiFHMzqIvFhRyGrpC4F5R0uzNozq9SCzbHgb1LGMYpBJBGAy10hG1qPFCYCheCXEpZvbCLH
jklMcAVj3R4W0OOcNLL2ayLkoYeia6evRY+4x0t+0K1JS1elusfBJy8jRQFXys1CvJxoKoYPEZMN
Kod3K+xkNnd/pYU1dgd7d5hBdcTYr8iSbXRefR+PJX3alOYYJ0NyCS8qx/HKQWJTylk2/YxUqLJb
x0EiCwVBsw4taNPZ7kDS++bpiExnmlw3ehED03leJh9zn8YRcFJ2yRRJBRLdZ/eadejM5I9XiqeX
3YoblF/cJxju/uG/R5gO8UDtO0H5j2QE7n8NSh/yZJ4HOJTcy+IRt/6gHzTu8Gsy87ajgG/Cj7AA
rFHpF9HLwKD0OskukixlNZjKhkwvQr2U2C/+g8/mLvkLDs1BymFHr0mpsZZ9m8WSZFGAgLVjl1y1
xW/8QUL9mx11+bK7MnI+EbBHeiDOS5VXSnRWzr9EJ8sZboolAi2NAn0h6FSPwZKWRPIxty1CwC2h
dVnnil94uALv9drJ0z/RJ6D66K0Zy6lWdrc9KOGfIxGanRB3hz31pVx0Zgd30i0yvbXSzro9Hh+F
4AuehAD9JD6cvDN0da9QwPiArLByKnQxz8DQyV3wgsz+9WeZ4tYB/hIlqXt7qQqNGIW36EuP7Uxw
L4CHAwFfCV0qj6FGxFNAbdEQFYSdLBz/fIsksXetEN7VfsIjV4ELCKyyv+IPVQpWXwUrN5/63H4X
HhQC2k6la8LOkjkscCregpMcMw8tCrni06AW87QA1Qf2iwYObmAYEM1JtV4SDPfYGjVp5W8DlmD7
imigsylFDmGE5NLRXzHTl+wHlG5BMUNRH72frnR8f9J2zNYjnpQDFqR52hkOBorrc013mLTijiy5
ErcKiZNl80x24Rj228JCLQDx3cXejWzxQ/15+SkPZWUomqN5IWiltst8z0VxmeL2/kIAYEyw80dh
53kiB+yW+gT1xycAnNE2iSHFORPZOVWope5YrNaB+Nxsc9G1TpMIxg41TxmAhK5kZb5HlMfyXwYd
Zy4Up2l3qm93c9yQtmqJcEG0QEwWRaawtSYlscOgGtiCA0QgeDojcDnLjvXzGenaFsLfp9rgA+OZ
xgciMPEkCtWYvCXEfb+U5ZJyGrRW5vMN0qxr7gQNarc4V3NF+k5zyKV106SYwL5e/YDYF+CQ5A6O
WPRzWm13VHbpZthoQwyRnlVxA1aUnH6xxU+DUjiepdjm5MXT+2vt2+do5I1XndsdCY9ttmNihuGH
ZP2yfVEX/OuafIoJNBMYDQvt4pXC9tyOK5KJkCBZG2bJ6GQSJ7KrWtr2UESufHE7g3gC8zsVGbtS
mUPfxGP3yQZQNiBuZ8VfXSxzhsuD6vjE0Oe9vspCIeelryA/Jz5s2yLGxSs8u9Bh4nmS+ZJczuwl
NEHUMRUQyn5ng1AbBYOD3xNhDTdShvSoHNmC7w+hF3DyzFVBXJs8vyU67Kl52zJRdhSUYx92hoJ+
5h2zOAGCmjufrUnIma+eKyzAOH2AQAySDxaOqbute6o8ef0/wVtKzlcppDcPOeAH/4FwR2qglTJh
38vEzHkzXQeeuDb8lrqXI82tOTRQ3C+rjy9S2IA45Tlm+ezBh04pW8lpftua0X0btFsvHAtReXh3
OhLnYZc2mXpWBjKaWCj/kur0KFJ0wawHiimEXRwR4jbnbWSN043E3I/r9SzfYsnboo+NmzrgmT4q
ewqsuRVI2h+97ZO+a2TnwAfZcjjtNXzCLFf81yHvqhWRAQLSBB9n6r4uqo4wGa157dDwKC9V8kcP
44Y34oFNRv5wA0NnTxhvZZyi6s8KjjmBuO9vYsMX6VuDTzBY54KxnYgG9IKPM/bL2zzZD3C4JvFl
VWwRU9TOI82FvEAidPZCWWHkHb6euByUNlp1FNwG2BnBj6Gq3VSUnsfDlI784s9r3ts1JUcqZqcY
wQD2kBZEXut4XtLtd8ivu1Pk4wbf6HPfnrnoPWDskRcpLZdWMg+dfphjWz2ebaBPb5o6gi7EgLnV
ve+4So0FGYG091lXAKO8itbKImlj9817kwVZSG3rhOhImUHKbJ6xaLEc3Q7r+RTciN3BLIP7/qOW
D2PbdDC2t9WEi7p3Ckx0mSjiASiWIoQi8ocZxDnklDgrU16ffr4mLnmPFu9q9CCu+Fre7MwAw8W1
1dQCBiiWGOkUX/ByI1hE/OIc34tem+l+DdhTBb/vnJlmrNQDISMma+enuoEo+BNMG9Z0FVBN3p6n
cYM7Dy/lJfpkpjIA7B9P6VWoAR4/LMIjEyJ9K7/RE6q5AGauXZG3DbyVUA/0fhppsTgDnFt0ulBq
FAM0xidyKXRdbF7i6kw6ZWta1aq4BOSOTckZb2rIH2jGtJ2f+NRsD58V+r6XLMigayjHnWe0s/Io
LLZAhgAPkTrEh4dPeA//Vv/KSgnHmzgGx6GFx13T9UIK6br+hXeyVyI7HhXIy12VE4+s4GI/MeMy
3wRocXNoolp6afarKRsqL0XAQStf8+eweHvGZ9M2+ZLEPP0DLgqdHBBgwymPByyWKbBvdMwzLUSy
Hkfo8F4trbSY1DW5gqcR30olvRhmd3hmo/FVAygR+Egvxg9B1xsPq2+FHjJeHULevwkErAb44o27
+lZy6UEbIUZyd0/UwkXxHg9l5vYSfCrBKiduRZ8pjyttxmiTBbj9NQ/OCweOC8CkOAH6AdIi3LW2
Ytw4HdqtIsAFcZTnWOeNpUP9+KbJuBw8eQ9puEj8dkXyY1il00B/lvbw/vOtFC1OQFYbRxm/wo53
Mbg4pNr0Krt3fXcWZek5I8BJnCyRSxda/Z6FsXO8x9EKn3uRo54jPJ596DRh8VwFCifHRtQeic69
3iq2K0pK8ynjSlIMjoj4GG7+eke8FtvyTS5ZlX+ORbYOzGeEf0pkPgUrbcfeDFsfX7OoYa1y9IRs
IjPpBQxweiG/qwjfZTQlITP4GP8uAzsJEzOiHWEShLHYBQDSzfdJ5b0ex/kT9bclikJZ+RZIMQ5j
0uPCjLtT4fzL8TQex2rm0kSwMhZIR5lGo+hNexrk6a+Sp0w900k/pcbQYIXXnCEFqHBrFkmpNv+A
tHPE2voor6wlRzlnVSdI4kRcpZuFav69DcyYn88e3r7CdIPUfpczcTNBZXeF6vAsfiqqb1pL5gMc
4K5Udce5dw3GhHTPuqzwb9XCZWr1zEHOV7Ed64VaIhEw5Jbhd+lekyzCOMCXCBr+71dekR6OSXnI
7E53VNUNoa2fwSXzh7tS8l+uMpVaZd0pafqomYWJTij/0zP6cYVZRttQ0ciBJi6Fr1zbl0qt0aOJ
8zoVRUcWK6HlWztfHSsJqgby8lbwKighOB4f3IXN95iyqXm7XH/Lb9JzcyM2IYcB6Q81NJLx+PO7
fIsQsCV6/BODa2lU/vax2iFD5ShJZ1r4/k1QA2dqV6pdzpWTXe+mhwEqCKQNqA8I+gZWW6WuL+ni
QcJbxlFmX0NxXHKXa/NWcDMlqhvst1cSciFFB7Gj8K9DAf78HktkSNlBNexKaVK4Sb9yBPYiF30H
758LCsut0jjgY5ksroscbsVLxrcwMGiNkIOwXNyhBcIDb2NKrXzBMQo5uPfXCFm4I6iUvfiSIBeg
mGnLsWobpReeLy4JmY1A8oae1MMOfu5IwMi8ljHLkIL9K24sB1fUlY0PAFoCSDVZTU5heFWNqfwH
QlxPXLCbpo4LQOKdqDT84Ws29B9RZq4/Zjf2NHLo3rfuC/w1qsAKDd4OA43+4UP/Qfr0DtVPD/5r
JRLzGjuObgHAJyOUc4Nz0N1Szj9EsNYY6EwGkB/g9xUgH80vkwPscINtMAtWaT9IXV6r0i6nse0r
gpl3bczp5fwRKrbx+loGCKvrn5VEMo6+kA5TarNozMDGKmFtjauaxbTnD2Ez1XqaWuPPK4dLJ0o6
Wm9UnT7Ob6LUywQ0cLE8I38mA8GSDDShPZ2KwmER9OcYca+HVMkocK0e41I8igVl5hsupVJMXTWx
bfB5zy0fakfhM+UCB+BBLmaxy7S3C+CRppp4LXpv/VVWsHff4VEA/lZkIoG/CZ4/XODmwmLfTN/g
3AhdkwfhnJ0M/G72gk2ESU4s+g90jKj1A+ez6FRzGgjd9shydkrEUh5U1lA7G5hJ25ho0SNtBv0s
Ws2Wsm+vxF3pcd5ihYgcsCN5W+4k9MoL4xI4pMRgutyttgnRHoo3Ypf8QOTh3mF3OgJTOtAEEOkZ
zdu+mSKeGWvdh5iWPa+b61fdJgCZ5Ty9P8WS/93hviAwwcgbLNILk5gsnH6Yi/YxttZ+WUNhSm3F
MUFijuVkz4/kBxtUoelyA7QZcnZIcdcfd8Cekhz3OqDCJfW2TdC9ptIxRWFnkdHcrTdkTRlRSkVV
HneUypLGgUolwfcQSOBUuKcvOFt3kC1yUROfa2ZI0u9TEPHE8xLWYQs5fXfIn3rZRYJDyOgQNCVJ
A3hxOyJz6u0ht3iXVrh9KyhPBbzR68wG+imJ/S9D48rqaBlMNZ5krxT+hQI/PtPHFHbrVtcmOA+R
QljEMTQntL48zjqXGdmLZ3puJmMPS3zdmOsakgE6LKebZ+7iA2AGzhBh55us4Sg1W9YfPlgX+WSt
5vCdkR6UDMUmJO6sPWmHNpG8Un5MTHqw86nNpziZvAP5uw4FrJ4dOsnNNUi+WkL2lvKZix90LilM
zmo7cJG9p5V/xGKthNHXb/GkynnSba13pl/gfSiZ7Rr7e4CDx0+rL22U1z9gJFd9spHFN2ASduN0
1lDGmDQ1I3On4dSGRqelEj23NQdSEOILAaYJQNtrHHUmXgKjvemQG3p911tkIGnqYfEy3C6cbu4O
xQX9V72K9KThD+THN0+pR15wu6G61XGkyl08byTJD0ursWWMv3wsSlPWjq8c7s673C2En/S82fKY
KHR7RiLc3YENK5C+bqOsd3XFaOzRyzpG1r/l8eOp69bZi8RZvSLElV+WJZPbTEdyDyZloquVCKJn
goLAZrTt8vYF3PbabWcWB7nifUhBhqf6LuSI6oE5WZOvqJdbEgTir0h8OywG3yq3Y5GSiIyLgIBq
5Lb09sUSViKbu5WlQnecUzQLXd1qU0RS+8xlEV34Tzt4fOXxM99Qmlv2RvLAVjfWfEimCaXrrWKf
c6jI2nKU/UzaaC8i8Yp27brEb6WCtNRLk2aE1gf9ZtveUsKtXJ8mPFzEW5jbe8e7r4FdgdrmIVOL
64EejRthSp3jkkfFnH/Ng2lr2hjtbueS/z1xlJ5Tr2fu0J2SEVMye51hulPmsycUQN4QjbMlRz5E
6gPYigkfnVN1/pRiGoJCZrLaopoC7ZNr/dWNwqonvTObZx+sHapMBvLqTmr5Uq0k+0tGe0WytUlH
DtZcAWA/I3V7WCBUNcWde5g/D5oq9KAtfKGRiOFYxEdDcRhNxMASA6UOkcxyGioIlwhhwRwITOqQ
uBgCA1ip+X8wlvLkaTGvFMm7PL5Gc8ymjIninnXXnGcpXrWWSBC7NFUCbVYTkh47en+yi64bKQ4r
iblN+/Ll7iyAvRGHHVS4cULatSGGSF4r/4gYFseDYf9KdVo6Kq4aQzzRZ8USp/gZQLABe+2Mgs8L
buvL8/SryEbhJeSkewy0jyYpmEzChEMHHOQOZDbPKWxrE0UirmJsL0bZN+2i4RmMCKXj5Yznaeka
89odPSoAIAnN2BgOeMQF6oqI4wIR+7G4Qaez7ocJT0XzA2+IijRm2Ed7W5qC6fQqnM2h9she8n8D
3/cedGzNUfvLTtuQ/Lm4uEM8xxoquFkKxXyXYeYqHTl+djXagzarCyX8VheWcURhWwn0VQClzvWO
Z/KZYsftFAzqQyJI8EgyMmjfIxfP8EXLLCH2ds/Uf6Ogkr9/Hy7Q+nis6nprpwyW+Y8Lpm7rRpaC
PoPex42b2f2NnuRIL3gi8RCVBpRXBEbzfPfDS/DDRyZW+Chsl4xoRnDkGiuqiGqlWO+8oeLi/Nb8
0Q2WhRi/y/mUUbOzY+HAuS0txwLkXJWr7JO0KFZz/VdH33PwjNkmWqgS113HuCFCMFx9Zsazjj0R
b6rGpdglzk0A6HTHGA2cUMX0pQVp12CJeUyiNhCxFEeDcRyGuc3XMwol3wYR//1ZRLd4S1EPoI10
HZGUVqXL1+Ep6/a5UC71gHci5jUUMJC6wCJ6CGzwecCu3c378xrttZhzhKtbMoZLgnZSOYjxCMD0
3Z7f+cf4ZzXR7nPet5cyMvmf6TOCxFOLchs/AZEFbTa20zyuKgG1dXkON8iwii0yR2tN8x433JSG
8rxDH8lwgzFMBURpHhPLuLSNeWIiSEdkZeLNYDsiYIauZKanvyZYpAeAjWwgMsQ7rLAx6ufxLYKR
uMHEbyWM0EJaUbe9dngmjGV81xW5K9Dg/S+g7q00vWV+admZQQV6Qge94c3M9HRnMjr/ZMq90iLt
uDgTblLSfgZIvPKWryZrUS8hwCnY1aZybLe+t5GJza9KZvuyfKcZHas6+xBPGQ7jj01VsWousg7o
YwB6yEtPkDcgW1qnipVibAaONmAy6VqsKL3C2xXt82YW9SHZRRwHZzP8ys1eRsmIoZ0QneaQ0wlH
mTWEP+YRBFDAVFvShUNotowezIED7RcR5lfyeiRlLXicfGevNSV5YfGJovEYWymRxXh5bzDhOFve
dQMVHTVSZiMzTUJheeezsYDTFGQ/Rw4YAgvrOG8iUXLZhYpsIrP7mOPhPqCVMfw9BkX7lYfTteyv
QdIzEtXKvYGjX0sIbv37atrIdTgmLe/1fuoxD4Sj/K/pVj7L/f2a6RfXfU/GZXeSQaXXFY91ouJp
gIZ9bZOm/MKucmGuhiQIocv1LB0y2EulmXtuSDulFdn85nyDW7gBfSm5SH7niSNohZzz1zwzlK3Z
fQY+nPjvsyngrTuGHfClt1hkvCHH2kvqXDsWtulC4DEMHUwRwEsmqsT/AYBJXCbPTTcnClhFTAci
9yOl4OD8LhHAOJi6SHFWLRTotjEsba3wNdqm4JJTCq6D+hk8zXyWX6xQkb0ydYcBhGK3Z1Euu0VL
l3JVeNt6BimRMGGa278p1Ew6z7FczmuKZ2YDdZA33M21lnRt6jayK5C9oRmqUeLi1VzYD/MxsvPP
h60CX3SJVyGGa4ER0+TYMjJNgPtSO/ECJOshVkYpXT4BkQEvvBCL5Xeh6G7hEhJ/s4Sah/OC85we
Fv7HF4dr0MuHBWZ/wkrhQ/1iqQS4ect4b6zTZrEOoxK7jclp5lK0oN+3JbaH+5x+sh3AWWv//rMr
R6r7yVlvFRQegfEkNkmXDxF6MwMZLpsFIeWfPCh4t5UrExn68Ft+bZUZTn15P9bE/IAgPa5odfHr
+pn0GJ4aT20wm1zlcb2Y+WSgp44oL2jDwQj6Xg+qFJ87WL8ZMXdiDsJrkwXZAPD4SpjzsfQER/Of
Igo1ZKnA1t1aFt9DcCyo3i32dvX58Ai8lBEdI2FwwimICqk+OPTw8jYMfJ1gdO2lfY6UIsfqJxiS
5+Hb+CrGJApUb3ILxb+iinXJfhXjzC7l1zmVMHq/zzsxH9erm870EXK+jqeIDwtD6msZFy+0bTpf
50y2wEcvtLM5Ft0qKAh8QNkPVBbmd7hhdBOmk6WJYvqRiXPfQCCBXf0EurBfaRysuAxKu5im6xdX
my6Tb2YWInXnAlIDajHp98yd/luueTxLZQEIN6QOV2Nn5jyFINO+gANk3WT0tPAcTfhUWwIWvL1/
bsxjzAtnLRamPBy3jyMDc22IWJ/n+W1CUUUkO2NGCWK314QP6qy716ZpooOrRUG8zcd4stxNxUEz
xVXLRRHgz3B9s7YuZmyKbNZyivFW040xI4jB+tU4J5lRq32d/ekkKMl3A8hCxyfo9AnNgH9cQsK8
ZKFyb6VqcR6C0BaRTbpP6u0asi/mPEuM6Dnhf7tnIzc/fGGgA9i3aWGHTkphyEnj8ILAHo0Tbenb
3XGVjjDQrIzbuiNDLCpZUAcf6G04PoxksT8S1aP6JAmguvspy9R7B/zXzhM8O5gmSv8DfYpDM2Ma
8s+VdHQypuAgE5H0jsYBfhvYVugsUd/y1iIAzwPEiRXQJKCSVBSNJKulDwhhDCu8MHOq2t6RAWwj
a7HKoRZVKSUN1T2TVb1ngzHPRPeoE9GDJOOF4RtJfEwBaAHGAAC1Jq1WuFepc07jDaZjkkXU97cr
LBa9so5gWwWvK213Fc3TB8FccixaZkHC8xB7lvtRaiw2CslZPq36fPuzlbkF/n7hSUk9dejo8y07
POGOemJ7T9egtcA/COjYEazX3D4ACKLZAQnoCpMmQJYDVWwfurIobmGgw8hDp+eWU+rhnNxhjy/I
s7brcutimldADZ4UAO8ZWSIDGIQYC7p95iVtuEIrSHYVNc9sEVj/EKIDCFi7BQkCdvZvbCkRx9hz
XgNm5aCKmdUYPky/SFUSL/tq6Nfwewkp+zOxgzU5iEm/9dHkEZBo3RbRwm1P/SwMFh7XXLNZkMzt
RSpeWvc0pg2TpWCnDlxIVIxYi6hEnJvxvt+OwaidOHRhO2zgn7WyRvo7CwbQ8hKCl5+jyPLB3UBv
dI1qAhvEth50LqPYSno1HQfZBBqhjLklSpqtJU8skN1grctb6MK/0bpZu6kGBDbQ+eBjS/bgh+H6
VGoQLao4y572aQfi0LZYTLn2lp9ZHbrlZsPM/a/N4TH1jtN3Ml6GXigFafc1/8rQ93g9A2xZ+JpH
EuxhdFb9O+0DJqhT/ecTloVBD7eyeSF4JTyOHzpShbkzwtJJxD37odi988vKMU8eWQE7nJZOb8k6
oSqhBo2Nz1v1/dwEkpgs41sAukzksLDSVqtV8HYiH+3qoE3tDpgjzn++fA1JsmCK8syAqdxd7qAR
cnzmvEA5wrG1YWCeqfW0KC8IOmaoqTpQEypiOPl3fp+fN1rmuM3MKs5HGNqGohsqhF6APVeeHPuq
8zg9Ri+eVEB8tK+4HUGrxq64zFFHfYNhHnFjXDYdnt51ljBUtRAUkRZBUbtKhSnjzot2joL4QSIQ
CiUedUoGr9Kaf2ShwlXDAPQr8eymcQPIw7AI34Z1yki/EJzbGbeLt7qJWPOPZxMNA35Y4c7MD21h
hOg/ifMe6C2u3jEQ8TFZ09gshI1LSZQnoj6eddlV7EB0qlZnEs4fm44VbPD6Am+RUtPFj7e1vdBL
GfR+fenWtxzmYHX2ZqtF6A4tDwRfm1xOpFhZXd+ThiskPQ3GMNvUD2g6dYnyqjnwf6BQ6jr6u9U9
OqAJuPPzJe9x+COe1NmG66WTGAcZL0HXk7++YTuSCpV8cAZntdVTcpYFN6LOp1tkJqsnaywEEwXx
KZvGR8chRnkCXFbRXy2S6T81uZeuj0XrpvL6i/7Ly9WWqo+3uhR4r0y0gVH2TxMV2B9sMCo5Zj2L
JXG3XjJBBparuvQdSX0qB2+TyQqCFTUVMkdpgKoILaWtRqNkWrIFJ6gII+eIT4PEW/0bAsy/e7uJ
WG+1vnk86Ff7po8azeKaNROr/GQMcsLVjSpMKmueJcDt58SLyrI5yVMGGpDDqSmBxa4JthyVRizw
kwWsE5OtpzxAFhg17msfwA7CtPUWpK5nQFZ96O1+RdMitWT1kLC+6zM4iVJViRItok8mq1KH6Pyi
hU3BFSwz0SEo7l80vAgE9EDEjGWaDvnYz60x6G+lOU1iJFmn8nu6fbISC4tj6dKFtncYhzPFrpjz
hQyM3IPrOmVG+oMMfauxQsBxaFQ5/Sb50Out7nuE9Hl2Eu6IGCoQdEiXaIPENyfSWAb9XrYetLoD
5DSLXo0T0hhhe8WrOwRR9lKbhFhW88fSiZ1YzPp4k1Hws/gVcWa2a/oWlP+bQa4vPlt1oWk2/PG1
/FpZl0XRvxeSrS/c+H0QrM22B847jxufxu+KDbSuJO+R7dxSX0oSB0wU/Whf5/uyNY8f8NGjsINd
iFq0iSF4UdmH+YH5HLQQW+5pnd39DN9C0bN+e77cu8g+gPstqB8qSWNZF++YkesZL5FPI1yCg+Be
GQD5tgfpjEMMhtc5kivgLDNhDgttsRqLPGVvB2mIN9Dh54cn8sBFKHgG+hTzp8X63JjmMqEtvWU7
fxEQiTi7cCwzkDR0PKo5+06YlIMTAT4nEpvO32nqdteEZRN0Mlow/D8ZMIhQfcIzdVEmLLXkpKiY
wD+43K7PwcYrQ2W+z4Pjp2zfTxZc4CMDsadAGOVDFa4sEG4URAr+VEq9y0kEbeXhukHkqcYynTMR
NfQXfrWZK9dIXHnGj3qjGzLZhAky0scJOYRExt5NZCY1mex+v7UZsDwAFyGlp21zpfWM/bzDZzPY
GrOsEuqjYvdLOEkFg9TfO286/vkeSdbz7E0g6vHunY0PjTz0lmXajQkY6dLr6WFqS31o85S42B/G
glU7KUA/Q22pgi4vXDS0cM5e/0YtrXQTU1VsSvPijfad+ZynPNiTV5iGzvWjEt7RQYBBBftRcMkf
+ISOHNvAsk0gSjyKDopqonDh7VjPMCyV5vVcuTlYiHRXnfZlt9b59D8vX/Ac/2ilaWNXD+vDYpZr
4hiyWQEtblVRTKtljsznK1ShzV/QnSjuttixsEGRp8zeT/GI7qllI9DFCCsq/NfbF+5vqZlEtlmP
0UNzC1JFGAU2UFDSiDz+WEjaBUZ3+DGK4xFyXaSIlziZMYGw7QFJ61WnUrXBFLsNAVZX1v3waVt6
Hu5FWdTBdzvM5wulw+IVnv4a1dGRx7RvUH9Y27S33n1MEs/EIOvTdn9gmS8eOZIXf9EQ7DPUBRi0
HMy0zdom/IW3c0n1dmVOAtpoooL4VaedChU3oYXoEVLDJrVV0t4lx9NBL7tCQ6rDWJMcOR2JabXd
GiqqmUUyxvWRRqRKf0Ef2h/fv9j+gwmL5mLMYZSmkqNb2rGvoNBbnmtU9iuu47Kxlko3dgZsPllK
7glM0wSdWpScHNAWbmjrOMv8RtHR4ApDxjMeSSuj5F7IsX23mRA8P/6QoHMfmzmOqEpFfGDg4GBm
ODGqwUD/g3nbSA7Yl4qKzgK+tgC/K8iXoo/YR0Bf+aSF5zh7ShXRbSEJItd+SUfBGPRSs/88+9I0
t4kecufAfr7sEpj4ndHYPvf9hduaKc+8eoug1BP5kpnSk09gKDqQWWBA7p6MfNq+XtX63YHZ0Oht
NICbyTrl94kOYQjYqXFiZFlVFXfwQXLvHtAcikW6Hhb4JnymU6OohzQl9/ubDukdTAdq2m3POSKJ
Bgnjgplt1xr1brhLIjYmBRvFoA1d156SP/G54hGUQLA0R4DZgnKYhSOV3Lj7C2x35uBDG86CONwk
1ERcEVX9zrSRS47FSpQd2MNoRWQz7Al69BU4pqtOKVuudHGuUqMI0ST6iwIKlPtBdrpM+rRNKOE3
gw5NH3h249Ulk+SJq7Hd3zq0b9NEOm/CVUTBQHbuArEWN1dI1MRSbooW0KDXNCe0f4l/sGGHEMcL
ZiTG648zs4ScpDiWZYSwhege7BsqTl30I/Ry2TIbHwpVQil/lJL16P+6QDTPv3CCpMjib0Bu1flX
Vmg4vobibl8SFrZ6RNI8iSiflmygdPzGDH2p8UJ5Z+WmX8d5Jvr+Uw+nitDtOdJqFTYTbsnn0ZHX
ACfBDFWPKJICED58zUepFEZItR0i+vrU32yHCPgwHwAMmeX9XUAUXOybXl6wvZwSYZi6HcJ1Usfl
e12OjhOpq5nX+S0wmCDSP+zo2E1DI+9Igu10GtUhiLB8YkS+RRurgpXk1Agzu3hbbCRIks+VyTHM
c+i5vS73o93vHZ2km/SlQwAfDK3U7y3Mo/reUoHy3TdsuWBy0taUctmRieHbfsFC+DBwH23SmbQ2
HVwfO77xaMn/8prPxCyO8uTGatzxRMZqQG4HL+PpszXl1kQcPcHJY0YXNfLDjFy5EsfgDDYxjQSH
pAbV0+IefnY4IgIqVPNDqPtN1YvZ9l9hSJPowS8lsoA4CpX5tfJzZQO4KVTDc+8nau25s6yW4OFS
BO9ummFRSlP/NF2ND9Gq1NTVLRaTCuF0hJyVQ0WHANQiSHg3UW1tXgOAq9wr4kjPGMjdbBumNuJK
VeQJdqGIXihL4+8SAPp9ZBeC1qNVZo8lV1rB2Yhmi8MCJ87/OKrJijXBfDdEBTBIeWTYJYQhhmSa
kpM1t+omHBoZAv+Mpm5jR/tv4U6+O/Q8Pz8dn5zL9sgp08CXX8Tx9zDs4sUhhQqJO/hBi/UIgCXa
aNSqe2zCgE2JGqvm+MTwjGk0cbdjRaEGV8U4qkc5f8xcxldGhMS8ditCFqfAWqeH0gSC91j1jp3b
0YPbfJOVFQUQFN+uGEP+MzWx5eLlZLp6W7sody9dHHcVA5sB1KrDCR5wlC+Ykzf31dWrmqnjtT3y
AO0hQRNPOAvW0Y8n4HeGYZzkBgDpjjIqPjnREZeubNu2Biw+FWdrpdvO0vu/NJLYYnODJmo4Osoc
Dnjl498WRE6sEh9gLLU1PnjNkSooI4DLJbEUPcwdmVRx0dZeDetLaCazJWBN5tkL2Do3AhIw6aXV
HliTG7gPvSVyvjKT919EjPt7bZnYSWnyM+gm8U0FYbLAd+YCPiA1MthWmZxxtpalnbXjTYDrNl/E
vHtvp8elTOIAsIhBUyXo4NeNfh5AAZIOyZEerPFtgJXFSgfc0It8EoTWAjpGAOi0pquwdWZ4E5Fd
fJV/x57VuT4KnF7JUGKMqzCl9XZZbICCRjMK9veo7BMZAyLNDc73QED22gXdOpsjA5rbXuQNC6gQ
9cxcylN2KDgY4R7yC4d/fR8RbMQFFrlEIA2KxeGJWHTP0uafD56/DfRWyN/7EqoQQrjwCds/970C
4pb+uRR1qGUwLiQpstfOgPiAbYhsqIMXX8rbPCQ4k8GlvLEEvYSsnSuPb00dVyFUSllUV9uhY3E9
Ijjw6ICtzMtk65da4GZBLpVVnzKAMi49PdIoaMxxAZTiqrE9ymgHQvmPjtYDfwJZWAL7NNDioFFR
rT8tMLLVqnYFhi4irpTRfVLA2TghoLvoKG3EC5p4WA3h1KOdrfykKkHMtvo9x5dg0ju+dwQgElUx
wT3AOLPjJJxp/x1anI7dp3sPm+FLw+kRq2Ub5truSX9SVl+2hFPWvWzhslUnkzSHrpkxUFk9FiaH
UbXXi/7+uNp2REGRaYOOm+LeCRK2wFnR0BTXLbm8eq5qOwT+kY6WsOD/XGYwTvQhG6V4wTl5Yhfi
Zrl+gpeNNGJbEmOTE9cYIcHUkzVNOZ2stgOhXG26qNnO2w/Wwltk4q8uNQix6IqxRlifxNUlRnEu
nYfBSNWcslD+N9G/OJQcmT8bF4Jjr/qw2VGWpea8bVtjVZ5obzOzb2AhFT8xfTWgDg9sTboL3fPE
rINhHO0N5SMe0YDZT0HVDlZoAglAewSYb8ico41x7intuwpBuezmspIa8C3/QSWRPKh9rewFsnlt
/IlTBUq+IQXX7i4BXoHfTSYkMYoUVSqKi3JETFndnetMCYbex1WTw7cl44m+x8aLqXlJkIgpxnVg
Dfqn+mmlRsck0Cp9V9E3gNmr+J9ohB/UDL/r+Qgsyt1DCa4Z9A1JZn5C42R7WS1cFXhMFyAbWrm3
Hkzfqvm9wS7tylK/9L7VPTcvdzoit3A8/hk68n9o32iRrYC/oXjeyDTrkqOTxt57epxUQPv/PSNB
lTpf4u4yDiEB/j6rqJ7/zckfv6jsoSCFeouShfYXVKbGcAs8FmRIFKGqb6HVmCKIm2mMHUDfuJ9m
pz2xZ73P/d8kal7om9O5+DsISGIH17wxUoNfNXj4S7t7mCgAEK3ReIM1nsQKvGPfW7hdU010d5S7
NDOT8P+bWtupavRetZKDd4UQb8F+2jwhyp+rDsvGW+m2lrUIF30dNIIzFx7JkrWobtZ5MhFLuzOU
0lb6nUsqn2Na5boT09tKndFmoHsi4GR0H+qcV8iOqvud7ZqUDTMuFHfDRbM7BWmZ/ZgEccnCksQZ
gqORB4HbnlndcakNRtuOQw2ZkBpGIHLNZZ0k6wfagdjHJWQEcTBqz/wuWklQOPTmq+YrpYznHv/4
Z5Wmapu/npojZYQ0QMmp8rLVkdYacOz35C+CYnHMKY5xf+ejagTFFB1HpRnqtlESC/P+e0n71B0p
X35+wXZqTviigRu3xTPHPcL8cRCeu0sRaSePhNapQeo4MsLx8HIMJZhnO/CFFWDCufvL+ggj+DJb
F1PlEwu9HIanr9G5scmgsUe90iuOAi61Dt5a1N2fDOsTSnvDIL9Z7V9On3+5Kbv9v7V+ZVqSVxEG
YJ7imDmncDgSXseEtyfWKvC8EXYS1AXIHQtGTS6Tn9kgX7CXxjnw9KWoltmwGMIqv7jymNsshb3Q
EYk1NbJhGwiVojx4fDLzwmWmaS7FzB8JBRr0sj0NqrTx6o+Dh5bSyJnO0vk6O5cVyiY2XiMB0yh6
cTakWNr/1Snhi69hknnr9Ma4+Ulhg3hAj29XvCLLpTh8TDw8fEv0rL8YnZqG1J7NOAQ3cf4pfCDY
madMCpWend+KH2+kzfAtb0nNbXhAU3nw4TPTk876b97k5ERF9B7ceWRNpn2Bj0sXvKARiYBrjaGb
5fryWveOYUrQfRUGSKYtH5yjYLJUPkno6zixMkfbJqBXiSm5T7HKHxb6eSjVrFeFwSZIGTe4mtOt
R1lkATdk9B5DFzt1Gxglj88KqjW/TOu4YAtFmp2daVllCKyr8st5v3jwnNV1vg/9jCs+Qm9W3uNX
0mCt7wUISsXJ+aGTeafTSlD05+7hCwMFsEE1Pt3FSWZSMQYIYFIT4kZvGbklXu247vVrzQSsCs6z
9DTMc2c7YkjOKrVeob/zxNSEmmtEtu9uLQBW06LRL5qOu/FEGuHgd+h8pjW7HOC6TuXhM65/1Yni
3kg34w6wuyjwPFdHOsRrj+KHHpF/801VgvlClO4gXt1bhgmbgPTw5jeyJHLZlPVpPNRdontgosMX
5YTbIwD+MJ/jm0C1vcArgexhSFIbzpmZv4pfbnWA/qBr+KwCcLx3At9Fdqp+0/lw5Tlwf2gIyHEC
0UhJ0UOwwGXcopk1ETBWig+bvFD5bXoV94XEmB3A6I4ah8zTBl3/b8IyPL4pRVrBPPKfBSdjt0Ku
nIKgfjbYS9EqBjIrX1Rp0OMCvE7f/VycTWiAgVsT8SdkLHR85nxcmEqtselOjKeN6RQJ3WeTggcA
I3+NDrU/0yE+GKxYGJqfIUbKF1rErKWGmW1s7SXU0lNb5Z3cH1IRQTawie4BPWRAqGte8H6GR4J+
TVQWyq/H6pmJ4Qyz/HHVYSKqZ0/gAurYKQfIgKW2263ue6jy0g6xkLlI4Ewhgw60fg+dTDilLUHl
iEzB01NX2t4GgeJuvalw/pxeYxPcaHmnPK//NHWuagUOWKvG1HjYizMys7ZA0IP7WdL53wPW/3CR
PIYRquUALmrA9bcJ4dH+qUT4hRYFi7zaqhqndPtgNC3FGDuaY/AqJQQFBc+6Qdj4KoVk9EU/X2EQ
tq1mxYd3/5Q6ERd4y0VjVolmRpWdoUEWmAv7FET+TjJ1wVzWxOZPCu14dTXV032vZ1y+Fiqh35hI
gaBId3MPMEaw+MehLxnxypjJTmUWkEz0oSJjyBZ8ZdexvYksgSa7vR4jXCeUwD5bzZWzv33JHA2x
mf46Rvv+jTtWAK/2nOhFa9UZPazGHO8zOnjC2VNguxES4f0SUTJXZsdbWuwNGHeTCnol/Ef3A13B
1QrEtKLo3EydpyNHV9OYpassKM/NahuO8Ph/bfGMrnp6ssjJvwtiZBeHkI7xoQ3Jq28q2tilXese
gxJBbeftlRIg/QfJhUOKuaxoUkIz6q0DHXALX/HHbtm6zaln/m54JdsONNWC7RtJqKQsv+vdW6Rx
xxVh/Y+RsTpBdiIUCvGoWijTPgRx26m/cKaYalcuot6GBXkgUE7CHX7AuKMHZ7qsoRJrmB3joUTL
pzp868404jF7uWlaFIrdG2HFkL5EavFjQ7UhNwTzMdNe622hqAlygkN/Qpq7YwgRfvIdX4EO/Wge
lWLyNdy1ior0IdnJvKvWFIgo7QST73FAp5Xn1p6bhms84R5W/2zHhdn26l0JYB2i6x6pj15QbOeJ
+u2/KxluP8TYui/b99Cgk8zN35i1eTX1E6mE0PdPF+bNhvWVprS1e/9c2S++4qDSf9kuVPum3lLv
+6+Yh6KRqYzxy9omZQZxq7uewjkgSQHRHZw1VLqJhOdde4Z7E9+JerZqlDYGXOr8yGKaCJp9KGSn
kYuPO53ilra5nn36xC2Dm8WvLLuZR8qTAIFYFKwED176/RLKoEAPxWBRs//TmpQwKZeIlv4OyzBj
MPfYdG2y+6ZKixrqnwl82Azk6YkZ3Hbxpx1ucTZ2dLIHEZxnQdsW4LEMaG/1uRRtwi4D+bmmOqut
PnRudbJojnf/hp4odNeRVHhsyZcfQz1fW3MWr+qixpjA+80bnk8zth+IDVHltpF18g3mlYHJfat7
V3jPXK9bso/NN4hZ/QKS+1adQ18k1MrdX9cJ+ZDdtrHyzT5Tq8mP/XShFS8A40M/xfq5P4Q2AOFR
Egs8Ss7etQrdDykE50h7UDBfmmvDfLOxUjd6Uhb7fQe6DHCLa0zts4TgLJWHrz7FMBXpSRqI44bf
WNXz9tuV6MI5BYzWHfndC3xWgq3x1k6jAfe2AgUIb+b482ZusvPqVO/YcSTOe81N3jPwiNE6Hqh3
GeHPoBKuufV6UHqPcQ+HCkhUQNXuUO7Mq6EQ5Cjx7QHXMAmw0FEcYtozIpXT85rZrRbxKxdtP8Ay
TyiM0tGdZYsLKir85wecMttgiG32TQUtudvB1PtXO4T84JIkNCpyaMk/miMux5kZuXbwhZpu4r9C
/plxoeF6lI9Tm0wA98KGG3/ZM/AE5UOTvnUdaY35NiUrGrYURd5Xagwq35l+x6N+tk5A3zVXMm9X
3OTa3eHoz/hEyBzUPvZnouo24Z5vWSuUjafyrikKOFWMBPSsVA8lRbOhJV9lof9XCfmuA4zw58Bc
i+ow4P9ZcqwI1Go5yea9e3HnBJv3nLbwLH0vv4O1XdmoOKm7DnujSuf8wy0Dq54dlXUw2YfcXmEW
EG9seVKwkhCRAK9VgnSp07u7rDQJyO3zRMkxGjrehdZq6WGc+yZfukx1sZvXnwDnimGpa9znk1qK
qPtJ8qHdKJyzDtfkTgle/GYuxs3XdX1SVpIiIYpxm/b4fSf+EHcwyL14VMgcF3jdj3ck2hQXsz5F
w1y3JGi3L553oBlFCs4Er9bcxXBbnGPX7dVUJw0XFdS3HdWBVE21FZH8gdkLMhDJZRDn36l9HHwV
X2RbyymKRTQEF5qeqTjRifNRlq9xn8hb+fCMjkmqTL6oawFhTg0RbrN+TcylvxdMSd1AYpTjCX5e
iymPXZdzhYDdH3JsRoQxDoyWJNi3j1Jc32Ywt8a2G1yuhYcSBUZkCY9xcVK80W2E+qEOtnTIV5Jk
nX5uTUDFUytC5t2MAih/XHgEBbwjeaC+nJb+yF0n2Cn/m2lRcKuEi6/lvT4b0izJIyiQgeoq/0PW
HmmYg66vGOtYS27YlrXa2SvtimuI44gMe2FkaQx84ImhRb2Mk9Ue6cAab0x8v5Yoo/ayjFZDY3z6
ocxN2zOs8NGIL7N1gxz/S5Fa2av7IDb2Qh57jHtp5fJvRAX81qPotdLUAbQviKz/XYEY0j0bsSDR
iTN9QoVy2WyydQJj6TdZ6lKJGbiADBR9RW22afiP9G/boeo9jqc2QCvESFfcfmxrekqfkhzEtXjt
dbkHZ0T/OQUZf4xudXryrff+Rqir+hWpOaOcbWSyxPjMHsEIdIAqJg264eqG+23uV72mECZF9+tF
LkdKEJRlswModmyR22g+tmKP7i8X6Ub5GgIHa3hEonbVdFDfRvAa9s+cT1VaLKGBz3MrY76z813J
skRXPQ4Ktogcfr4qpGhwhfvg8vC5ZhMx5sN7pCNcywRxRzWziuzDEe2ku3rJpcH6MAiNe3M8BjcM
L3s0wG17tHaWBYxJQVcwxk5EtXmtoU4IAV/fszyRmFSLrRJ+PDSnP8RL/9ifwL77XtrwnzqfjcMj
3HNwhvbkapNkgftAZhFewotExEd/SdYnc6MfP0zCwSJDa7Uxj6s42us94vx0mSt6g5zFemByvQHG
U2juaAmcsl0gjkbMRzML1JBO0bM2JjItE+Dh2bHQEMFc1riHZLpioYOoit/2j8YwzpmgMy9KJaDy
BcZpizbpDhEE90ec6GWVuD/NuMu6BpkURjMwGY58zUIB5kr+1dWteLOllntrNKf7wo2AFroB74aA
0odfYy/26z6T8HRRj98lbyZ74dgWDB7npySSjD7lMiOIZnzrUoHdmQml/OoMcRx/wsUFWiJUNbhS
ny+lb345cIGvay958UUWk19RkgohHnN5WUyNN4K7LuuWC5itimhMzk5f0vpU9puRD9jntFGp7l7Z
gMmsOdn3tdn93qhE7Qxjaz/XcX6AtGfFMToz69eyR7QfRbRF6We70jshzEf8IBHla07WFe8PcPqP
9vFYK9BTV4dqpnTpE2gCWNXOz/SvQrdtjaLDWyiGdD/EBlYEa0LwSApDfggjaVCG3WIAawvq4mOZ
pZqEHcLk5VI/RfncKy8TyofKrNxOCSKQQYkOPZ7jGrXAVma4k3r505t+hydqloQpIifFH0B8/lMw
/pTItmQK3O16IdG4vQYqfZPYTJQnK774Y+n+ykMfCcgICrPrjgU/6qOMl2C4JBsyc6uGqJkKfVo7
b+z+woYVnv0gXflxFlugR6gwlcsJ7QF+8/EkeWzGCIJAODAOoA20H9aqE1EOduH/pqpNhwRNFfQB
12OV6TgJiGX5hyziCghyI/6mK0hGnE0452Pz2fRQipQ9HE7QPqqXg4GRAZGlhxXNYQYffRTnCjlg
NrxzYwNF+b2L43YvJGZNKf4PDcUVmRVvla7Zaz3s4FBtvXmNkS0ro21LZXiq6yjeyFtjdBP1XQou
tg4/A4UCCEtBEGR4wqmn/3pvft5YtabUXXGi2BgySAIzoF+MxKwRUCkWplSkCA9FPkyv5RKeiSBq
QRAymBps0izQKxZ8iKQXOm9vo2xxEcrGKz0fsZ/2l+kUWzQmANwNTnU91z6wvm86BPWhZcLnZxKi
g9yZkp8EB6y7CJGz4mr5o5pAXOf1QCWnooiZzQQdkoriZK1Kio3k9kWAgfTDc+4t0vQTkF/n85WV
rYZ4eGv92qhyl7ErzPRl9a9QtD57Ari8q1Wwf8RxadyB/ev9JGmZWBlB3X9aGRs8EkQFwttudh6o
JVcrQvQ4Bm8aoCcMZIgKbXWoddLnW0q8UtoEJ1H/T9A0is3BmVsy0yrQfOVpb7gFqRZ6j+x/8Dd/
/4bI504kjd7KpGwwK7PJlu1El/PXPQ5PN2giyggHrjdqzIKQAsaST+eI4xBJyskECu5KICXLrfmI
+1eBplhPz7V00lz5rR4yGhG91VCV1rhDqJil/tYXb3tm90BmKs8Aw/2U0FAkTNib276acHHwHfQb
2foTQccAq8M2VLo4oIGVNod7GAt/ehfuQAg1n7rllIbo4O0sK4q6Ohtg8/TZ8vDhbS4xwNtlxYQx
6+1U0Bi/jX75DQNEt+fo4beEHgS+KQFFO+oH/Tp7STWoz8yFiQpc7aEOVf8dd1NDGmqFa4dExzq1
inY0Jmu+hHYQ7uqInWo0L44VDzt8YhzA0A6XD2izx8XgtRaPv8swePm1D2cWzzZckXwBk3xZpP7b
rvQgAKNV1F4EBn33S9+6opviX7O9D+TE6xLhMx2moc3xY1iZTpy1mm7Twq2CGZQoXsBDKCoPy6XQ
Dm4VwM9ivCjOGO+CZRQdbCzP8LPj5/rK3MGrHtFjK8OtGgffJf1juTXyBjyuQsLWhz8+f8Yylg5P
IQk92++PHQRdglM8q5lCv82NS/rFv3gFiPM70f0zLg7in7A5JjtteVE95ilDHUr9Uo36K2AnJ/we
JuBI/cNQVARd6Cj9crUh3o9V+pW5m4WPTbCN/nxKiHLtMp49sUK7aDmQBeIzS64PX2QoGbt59ZxY
NarsVqYxQMMYu/v+r8CTAGftUT4tYjY/itCkULtQbVpyEw2PfLpRzc+YY3IlU1SNOv2ttxglKHdj
j3HuPe7Y93IO94mwrycjqQW8xyH7c1bA6/+RIaz1B7ujKPoupXw14F6Pc169pRK5ZdqKpIzrTCx7
0rhKf8hyWjyoe76pqr6ya8ABiSwCkdZ/CV7AVCR4gLzxyyXYV1qcSZtnD6YkZgUc8SjDTNKEhDDB
mOdGN7Yklp8qreANT/a9KM8+0R3Lojhp//tixVjHS1HqeU9l8A/qU/ijSNcn0RUK/Ho+c8FGhLof
aoFqOxe++A8+h917hFQsTLuBXKAiutKsuRxK2yK/Uzg0u/otYQ2k/FfdsJtW30mXfIV5zQhWpqEf
kUUx/U77xK016Utunp7n5jEJgpz+S+HUo7ILUj6qqmekRik6D5lofDh+i/quScFttXjdbSIdDn8r
A/Q5Y25x1pJiXNhfKNF6BhjBN9xW3r5bdkdR2CHruZa6WmKnYLyiXtpiNTPJSS/lunVzFMRG32b1
GxDSwwp084ToHWsmbHEOixOX7Lji61uscZW4JcNzjWapIOd6LfLJAhdNFCUM9omhGH9/D9E2BgDa
eN5MhvgC9hLHDQ+A+ygm2Dq99lx5IUAHWYi6pkzk2EwusaySCTRIIve8qQpKfJENfh6kvxfgBUYA
SCX1aa1gIDoEmkKpR8i//JxPBos/A6/oRus8jRQdQx1Dc9wmVvIr+kTBe5NooL2+HQft6VjUV/Cd
KdbScDePtCCsKuac0TNB8xuY/vW2RfMS4OzCdhjBeQCEIVu830bpWtBUAYnltFarqG0h6zYD/dJ0
RCbUVMrILTT3mncMJONY78EWi3fi8f4N0aYpzYcyx8E5T+okJBZaQjyeglrO+MusTzg0EvldXtVZ
3Ptc6JlPsExoM7dQ2bsnVniSMUELmVIPBo8RpX0MQjQX5Mmx0mo+9xUUF2Vyv9RgscACFhNFcVfF
xJc6T17zbiEIGK0tg+4+GWFgvz6Ym9NJ5sALgG35HvRdiskBY37Y3LLSEJnUS31u7uNo3zCMDHdT
a6n0uAjfmLovBnhGyxCA3vODaDc/NWTpvApItdZsnFRey7a6xCu52kaib96lJkL5F1sJiAbSxzy/
uiehtIRHOUBha0NVImPZ834dL0uTsNBWRRm8W67G+YfIITGgfWU/kSrPwhTFc1DwFn6l/RvYYR7p
ioiWEtmBSwB6zwfELzuippOTqYim1bEpO0NL+f/F6J4vIUXishLSmkAQUSh2ppLSI0lUCmCg1jVT
wsGP5cLkezY1lnZim24KWxMi7o1RO6E2biI12QVLZiuq6yar6oZ1EnxoRGsV8Jp6YJ4mc5NmCkt1
EAhnl/sRxoXTLpDuN1GhRnIHYJB6wQySdIsWYsCeMvXjaWIdtUKL+pm6j5JFehKjKamLA3a8lXZQ
QDM4JghDl/sUoPZi1FH/GWoPQuFd6noysWjL5pGRTgXXHh0kg29wOJESeoA4GyvZAl7ZwyCFoLuP
pOW1akmX5rzhElTqRU7NvJ0goX8widsyKzrv5mmBACoh9gFokga+KOn3Elaq2wsVywcmrQPnyrCf
wD+nTDnhpM7zB5PVQzfURJ6PJR47fb89pnSHxeU3TGEhRelTsrqDHrNjxPOeLSUJq0l0HOi3pz+/
Rr7W2X/yG88lCIzDNSCg6VBnC98xzADlqAn3r/L5gZ5NTLmIL9ShGYa46MPHNdMUVJnIxIDq3OqR
0A7YrAFd4JCZGDRGpx2gEQTvh65XChWSjQSMul4HXCk2E+DWBta96z2WWwMAEJHml6COJI1IauEE
3pk5WoxTzGVZs0x999l6BGL0cdgIrgkg+x9L2eKIq6D8KsgqkOHoXPTuiWBtCafnYEqqaa9U4CNI
YMmXgmK7p4JhhkFwcIsv/qTmCE3Kd1YLyZdlqMOd04hdWYbTtUMXQjihQ7A2fHaJMITbxAXY1UVo
0C7nj1sOwHAfEbrmrjqVM2Bb95qAOMNECoOovkyBPUVQ4ztax4PuI4kepWeh2rPUECrPzt0WtPwi
ahI1uuhu0QrI6QKap4FP0wFFdIetPdIDL1Fhw/RBxusJ253kJDQveS2CnC5K7IX/luOgzGylv0Om
tHfLz+1XhYFhlIKpEQLjhOTzJ2p+vtfiMvznzLi3e/wQ+pG7+XEPFQ641jFiWlR1F73Bx3fEEhX6
XSAsg4kFPYVZypH7VeeHmaZWPDPx4psL9ny9rdj3k4oqapUEo8U2W+kMHRt64JcZpBf3JsmOrzvE
GrmExkpgMDSGasInNiFQtzeyfTIWDXNF9SQGuij6H/utLpC7xEliFCE0Ubs/V/OJeRQmr3C7aMzp
ubb778nSJXICyUXSJ3PDYBDVYTT0Sj1+Xr1+ObNoigZVntn/MzFTJEmjnKi53URXc98qFojj9B+5
NxP93Me1+I10AMIx88qFYw4RULJSZW+7QGRX/L7hDbYLrxA8k3SMQ7v3NB7brEQs798OoqbHgIhj
dmcLVmHGFGkI5seCwsQwXorsQ0tZ7nJdjkZX11NzkTK6Nfu2I/gUM8gXHa69LcBSGMZXZbkClEkT
9pj7cUOBcKlEjmOThfxaBGWqMbFytg767DrYasQydRBtv9pApulo2yVrptchyGOjkIIWE+S77Js5
jOsuosP17mflffEHqD/BHdTi5mHxET/8Z1G+AGTyUdPRTX+DrKQ9Y6fi7p4UX41mTec48ksLdtJZ
eIf1OTPdBpLlVTHN+xc2CrDVHtEPQvgzStTULdOWMPZtG/i/XIIBZ1Ylrr3hHbM6YSPF6PUyPXgC
tZXaveocpl7PBxZiigqeq6V48s7Y8g6AaYa5z9hACxR4uDD0G8CiFKhHfgXI5xr1I4yJtU7jx0x2
kyUbd9liVVp1Viwpj19PI9kgXEzCjOKbcBTqy6PdspjcZkCt4XjFuu3nfdCKk89FAQMZhs4DO4/q
lpZlZOhLgqVTX1Zi4XIdBm8i9R1LYXxe8lh0U6pgFzwMCZJQ8jfpfdcSaLWCP+tXl0goDvna0Sg2
e1cCV3M2SYqzMMAMVwmBVOIHp72eSN0OMEGm6sLlnezIcVAubNmGj3VIp6pE7KeOcKVhIqP6lTcm
U0/3PXwwa73akGg979ChOieMNv0PH2b7Bhvow52QkFs+NtuYk/bh/f2F9TGhd3DLHwvUCCppuSEr
BtbWgYGdBjUfxBzGzi5YxfaKPTwjptfe6mbjRyPxMOlBiBfWYSOE4tMOHUwAQ0zlHIdyn87jzu6W
QVX8Dhx5K1WlKG8T7UN6tfdYiSq9GS9x2HXS0L4xr5Jv2sS4TOqoqRoc4AatoT3oUnArhY01JE75
9r5CnbOw8JJMbGO0sKu/eE1z36AWmLAbDjK+2nihu5LmaO+TEbuRBghJANvnfPwXQDOPyuemIp5j
kN3zMblU8p3Hn0DqpnJjkjuJheAZSjvaAnCyHRx1ogd/BfYdOLTUryCzmI9wsD4ZfvKKVQp9QnWr
MJOAfrxMAO8vz6cTAI9VI+fI855BL+YRHNoWraDT8uq4CcB9sqceMxaDcBJm2SomgV6Fsx8PNuY3
NjV7QyHJeCyIkgHpoaU2WJBn5n/FlcCUcOg3kab3KytO61olAdcJiumtWEH8OlA7dbldDQt/HERR
1VuIYFg0btddlBF7eev+IWJN4PjiLZIMmyUNsrx3m1LpLUfuuRpvQLEoqFpR0ufpoFsmBUVHkBvV
+Uw/ZOtDbw3FKjQPIWJIPbKzMwP5YzQTQh+fQtSVD+vZR+DbVdcwVvLrEq8aaqBCsxw3Qx+PzIFK
HCi3za8N3FN6XCnjQGGM3hMeNJVCyx69+noqL/7YD7eIY/VXSNvqyndgtzhr0DcaE/TxEHADSvA8
NS36vjKaUIkcsRQABa32K80jivo8yXmXO3zpZLbPS0cCjwVAXLkBVIQFNqBIidexhJfsIDg9OOwC
SaieTSj3WN5eS23xVUDYzQPrJrnLhQzYhDtUrJfcygOKOAur2OJjwjtvWLqMP3LHelKQCPb63b/H
Y1Z+UkPGzFd1BKD7JHpm70uUODkr6Mu1/E/vsrgRB8gQZzSkTanvO47sy3fwwn9ql7UwsgggTd2Q
DmXzX9RNWns0GnKVd2isZnLFiQr7xykYERDMfADRkdtn4isshAi14WJz890y/Jew8V/rWniANPbU
myypF+Y5kCRL7/PTZe5vIDPAHGEHJUZM7fIiWsUWcggW45jYKKm+8zhi/Ei6sHPwkMpWfxxCjA3C
b3JUXFfTbClps4Roet0ueJCfeY0lcNAdmwG6wQpobnBNLTAxLCHTzRO0J2maPkXDOBJ1qfISLeel
guXj5p/Ekr+owPHEzS+0d+1akFdmgNs4za2LwPohMeQUizI+1tAVzTS33qF6TtnsnBV/qHR3sqfN
12wyvDPOXYfrzuI7aNUWGhuDk8u4Gl9HDGcRjVRvm/+a3DSQZAlXYlB4doMu5tfh5ODlZE/PPjgm
53M3OamACdOes5tW6BMlFhIuMcv3weaq3WKwjU6b3R5z18OMgWapCDJkPRwSJkzI0jcbq0YXnVLm
ZYy+wqUJlbOsaGkd5R7l7Rdu6P/JACHFD9tqqzF1BNJ7lpccEJ88ed/D7EhO3+6BAHrbpEQ6CF6Z
YN3wAdJZH2qgMiyUs8ooQi6c9vsSX0ixTpbQIfAp7nNXeAOlNb1q62XttTB85YRlPrurWjYnt1O+
xS72heBki2qUChYjTQI+o4z9LaEdNNEhJMen+5w0RQ6Hpehi7A7zWpCcXQiX6G8zKKtrxlJLyUA9
UsbJzrmoGEMOpCwOnv5F5FXSBVxfMYXhtWkPuB/aREjC7qaB1SdIU4z4QO+fJl/JrgevIr/ZEtA4
5i+HhU6wDVbqfCKMvoYNiqlCRWEHDykAUOEYaAn2hqGYMeDXHK/KewLzQEf0Xs/Z6Jl8GI9TfJvI
5SaDUXcSU2m1NMIg8LVqnSrywZUV06KQwpT/fZSlNNmHrUBoLhuuVfslCEKXnGOq+JS3elFBp039
KVlcZIvQglch3/Fqa83rbWUCSRJ96N1BTUaN+feTrUcfFJKd64q963IJ6Aq2xPdFT1+G4/ZIkNUR
arRQdposS737WKRdxCURHSkoLnNgnik8K9z4npMNgFt1j6w9w/x4iPoYcUgX8mWBtw9KZmj4VBVn
7dTDWHqrt/ICBZVVeDdW4QBbL0QBj3wnsDF8Ad7KROsBgTwwvZIIT3H281kI5MnFO8tgh+/3gftK
Hm2eW6jENb3MRcokBHqu5Ezesmd+M/gCHYxjRYhaOzTFTIOYoaWT46pjuaY/o25HD+blUubwDI6l
UWC/vEEKo3IthK2veKpRy1gqhRQ3JrRvmV+GZicNw+5hQaCu2N9Er75/MpqfIJWrwWaLcQLrS0rR
p711aoJtONG1u2nlyTvjbSphBHDB0QBBplEbEEGHhWkdC29hFbVnsisfkWBr8gcrFnNmSiIBxFMF
i0BxtyAG+Mz3qx+lT09wrPS/oy6JdQiGwTrSum8pjfSkfmwhffCEzOV7Uhvvnl2l4YpBsm0Kb4Qf
ak5P2Qhx30W0spsPh/+3QoVO77uSkW1SIZLAODt8EtIBjrNQ4f/zoVXVJqk9TTAovJe7sSzch3Ce
oK6fA6xXHpRfSzWOzCgZlGNlWaX9IrHOo1Lla3XKRjUYEMPDx5g1zNWiRRaaYLclWiD0v0v6kAgt
iEwJ9o3hqgI2fbQMpCheSuK3/Cr8VZ3K21K50+E9CQEaHOrnYKtFESiWAT2iYLzQKW+VvjdyPiPU
VFrivExo61rYi5grP73xPomIwzk4ZTVAhg/SpCyVrbBtKQ4VGpn4VgLtgKV7J/DqTaa9yIpvRH6n
cXiJXtkjPQiHdKaFqTaGDbyLArmqKIpcgK+b5iNrVX0Wj4FfmphNlbtKW7DDX4U6DSzHWjLHt9Mi
ygikITLKoEDxz2K5yZCvKawOhiRFFzosAxaQAqdDSccZtLGYEbsxyGbHa6ZotAVLs5wRFImRlJte
Zqecm5N1zSoMnxooI9b6phWASZrdv9UCWC6VjwWem9p5kyq/3o61pn7Ijq7BARPz3mgYqE4S88Wk
tNHkMQEwkfDQzJynAhL1K77/ZaGqOOJgLW89Gexmsww2dcWlcYruI2dX1pGch609QBV5G59UrNQI
+HIpU4YWmVyA/uQCSuMfcui64t0c7NNCEBoeN1O67jie0Jb6PcmvEK21ULfbyAE+ZLoXwIg+eC2A
uCAhlPl4j75OsvFW+MyCgmMZrTwGTCeQXhVnuDYmKd8FWfGCta1GCpZ//ILp37ZSRpr7T7bfJ3al
j/UflCkzCDvA1k6rO0r68f193SqNrrEdZHiHb1E33khy5guRXcRts5yDIyedmlfP9chWebfUtsAU
HeWdVAxf/5scRiamEnwqEXinVVAnuL9VyX0zRq8oS6+2ztppeVx6UFYVIydqCQYnVFN0KKoo7VDp
4C1z4FPpPN7bxsz270XuI1LE8h/hCkuf9u7CoeYUrp6+HYkMz+6e9lFN3ImolhflO2b/lHG7Fr95
ap+4GWoZo50Bd/xKN7A8i1TlGfF+CUQHxmQ2TQylLpWZado6KVfJIwUbtRsaZJOj6+4XMB/RRxot
VG4YjZ6sE4wiJhQ3UpS8A69QxdKEV6dC78tSuDbEmhPQr2QA18SceCXuwDL7JGOP5rTy0q/mtWPK
c5kn6GvM6gBfgyHo2tQSOk/9/p4OTz+CRrxFExigvjnmyjham3YZCjYvWuKT5B0mH//ID+ahZ41F
9UG5vVRgLBn0SDMBwxtwbDzZmJH84YmiTjGNdR3TLklGRfomzQ4I43iWKmCIzI0oE0R8zRjW+HRv
QtQYNT7PI1/VrjGZ0KbcuV8RcomtDDcmHrmBe2kB62953Hs+ClHf7dgob/3xr594+vDJ/CmLRbop
N7ES1KdV8G+e78RlwIxfl9B6IkBTxqCJjlTI5yytZqIMMJ5caNeao+q+aim/a93W/LRLmWj/ha4M
bk7GEE7HEN7z8UowU8xmgPK95DwOx2FCW/OiqrOnKr0GACkI3r0vo72CGc2x/MDfly1mmDrgOqdr
zJcUpKYoJdTkYlJxEn5KvTJ+8CGXaQg0us+20QTZ1YaAwrwcFQiyvJ+N7JSPGscCuaM9VUFZ9B35
lBPHklCHCtx18AywVMmuzq1RHBEHIift3PQQZf8+GaIcvgCoAwkjP5Znxy19TWME963dAliWHAHD
I33/5PCjUR/5mi118w4FNSL5To9NCcEZJRis/LIoREtMI4008DnwCUQCaTjvSIDY69N3IAyUoDe+
jrWdSt6SSK6H/kubxb3sKeiAArZllalreImqtUAxm79ylzroFc8N//qmI8QEN6ScBwBc/+J8Oq+9
OOWftzaUp+wCkVMVHpfhBv0gg2Ev0+/PvQpiiv/a6/XUikhOAITVXPPYe1saZewvibg3gJlY3cMo
ObnqXZy6Vv0iSQklpyIxXGvcQ9y4GAZbpLS2+L09nXXIB9JyWl1nIz5GMWrTwSmg/EIClJVIYRxp
SENraW5VmneMSvVSRaoed2VqFDgBbGdu6PQZuVlL29e8C2lVzDKAI2Ujh8qOYJc+CpmCiL21SXys
MDeJpIvoqQq1qQi2La3ZlHPrN/Zaom76dSQiqJXHYPqQVodGyREsCRQPxpMLWGDrTQdJDSEfImcp
T55o1O8IeiJ4F/Fn++hHtRFn9zXOVr1lMi+ttNAFHrf2NTirLIvxaC9aR4xu1sSXs/kBHSd3asQ8
BI8n04Q6vdo+nzb3PwstJ2f8Vbecli19AxfyulBlOtQLFM5L8a2gCPO3cuqve7Om870s+RSglnin
q1KqyOacFDPojkrFUSLsmWZ42veX6Mz8rPiHKORPflVV4g2AoKHSovYAUeeBOECY43Lw/KM1Z+qO
7wAfOjrh17JYACglDvtvMrJxlQ77nmpBuG4Xvr2ipuBHdZJM0Z4rhc2HgGjdTVHVtNls0hz+RqVI
Sq4uIjpEr6iQEICkFJ9YTdRiELeYJHBiBUlVrblybekoES/z0ifQMnqaeT1Cf7/gxYGPwJFQDsL9
JDkwVHo1zooXnbFaIre4+92aL1qOJpEEEbtQajfjTyOM3Z5i04TIYTm9fAEM2ZvkvT36E5EZs2yF
y/Y0m4T4/Y7ssLl+6pmxgUFFnIfI9oC8H/1Q+FbNYZ955KBtIuppoyDVTo6gYcBGDdLYk5Mkohih
26y5cylKXHGkqBgIi9uCKSPIwL4CNdExMwkCfN99PBKBKFzKW3hGHSSSGz2Ms4d0JlbrShdm+Q6W
IPtQXDYhxcfj1gDGPn8A2A8J61+4P4jIx6jwzGRM/SRMdBtqaVM3i1p7Nrvd/TV6dUHFBCBTuufd
kf9HXuO39MYuEm7qqOfbn5kCydvTxN3fmfi/ZjUOxZskdMCWYuGGcL0TfF903tpimllfC2AzvDWx
D0svE91iHpnuPg/EPSE3xnunlvxNbU9Gqvhg4oXK3WrtGlQSI0QScVGSm2Srx+nPVLSKo04iNpSV
//guitIJDvPpK/oo/aCGuHt4Ij8Gzr/uTkqFYRFvU+q+PedULObzKqvmI60kSHBRpuLTDgEMnJIG
B2VcxxayJiygF70HnzI1XFPeTU9KYqvEmIpQ5Rd44b2phBgzYeRKGEvdl+Ar9fOqFkHuPrsuOAO/
8OYpE3HMTGuvJ/GOrNglAqHSA8EyN/2EawlFBheg3Vo/sTeazrMCZAURbuxh6NyeMuV+gi27IuAL
hkVGX1qApDjrvpcqmS+YVKuyT9H/OYZBEniKJ0ogD7MPGGAFCfHxLNkUNijqlsfTKzSDEjWsQXDH
g+73zELiETlIG8BcXgrkz4+x0oj9uV1jkt0XhVgeFwb9IpFp8Pm8ijeIdvS15UIG9HR8uOkR6pgO
HD85gwnV+6rVVhTV+KEj79s3RWgmeAZZm0Gz2CNUVGc6XAoAJPuF1LJ/2EZiZ57eIxqXcM/H8ig1
Q2Of1Cc+l1snvjA6zPtcl1CJ6WZt8jLtWWX5LAQMdNRkgKxYpKehc0jw1IPxMhZqzSdg0Wl0OaTi
upX9uygcs4Pgwo7sVe59bewqZLRgRGYetniBOOIiNb1wviQjJmgWpPDZ8GGwjEEniNT6Ozncbypy
6+rYzP7U5/V0dLp6FszfdK3WhiPYv0QgurSN0yh5+hk57KJ1vZnSml1U/Zva1YQhMLO9dGcfGRdm
wBWgN71PqDhyKSSpUake0AJHaMJLlwTQcaebPla9MvW3g/TgS0bGqJ559s2LYJRGes9MkXWQ2gqf
zcGyZyedR1Ut0YTnDed8zFf51KyG2IaiZYZUnAO2XHAh8caUfKsYG7Pvu/ntmyAIeDcVRVFtuowe
4wZEAkR3dRcZq18Jgmsd02QWBZLmwyYuzpOFrJmy37PaOz0BwMaUUdRUQnlqh6ov38lIqBOwfEdT
zwwASkLl7CmTdQuQC+XeH1XljqJQpNNYl4csxdvMxMRgokuNLKtQf/2srPIDOVnp5gsDTo3zXpYZ
wezGOehrMpERPQYF+HZmhr45C5kvRxjDoRbclMFTombBLwoA0kcnvrLYE/P5w5jPMYP6CbBiSJyC
Al7RhqfeLvw1HeV2K9ZmRWIVGcmfd23nZALcEc1Spy7h+lSbPk1b9WfLqZisqnruKXFI3uwz76FM
QQpsvjCoKwlPWqwF9gd+VEF6li9XEtlxbmAA477Geq069bXjQ+rFdjkoRikJlA2+LXZu0jOIKhT5
f1Hh4g6oRUSWLPdsqv6pdpQW0pzvVY/79vKijNOBMc3DFOSuO5eGrzAmI+ZuYL1eCt12ecnDrOLK
7KU+QmcRL2LfnThOgPPgQvr0jtSTX2VN3bASA+0d4lAMMW/r0fZS90x90IO0+qybB7KXP2Wkr/xy
b7KAIDMDE3XzgVyV5cl46vA36ICp6s521OHS/RaVkmdcXLqP2wwpJyZ1leFtvXgnI7OfovVSPXnl
T6lB4dYevRjxXeepY/kPI6P3mtM+y0E6xCNnWT2GeuCpcrxZb6HI1F/F/v2J+FlPTPaqkuV5XjHB
lUkdkMqgg3tazSsEEqF3AItuMSDQS0ZGC//moXBU1iB+H//iW79v9Svfj5dxMOiLkaNG2H8oPpYg
svtJhcL07lQABcahZQl8vDQbQoYWfgyxz46Ws6dM8FxkGClV8+8uVp176MR4tdKFMxo43RvEkqPq
zujS7sGRZjQx4BkUFe3O7j0DC+sMfWULXjyiKBKHh4mc7iLqbhMXm7uqsg57IYHRkkXDiJXQ/aC+
DAMhY6tiOWparx5KS2ONfboQxsOoeSBM8MB/FC4O8K9dTyS4UjxCWeHBnvRytS6VS2BX3NWaGR6d
P8A+V3RfY5oymKu59DwwZxZXW+TBB87Vk3lb3gjT8gI9G4yM6ccIdvYYlSwFutg3xwoNhzO1tFZB
dLXjpzFT+lUKL/z/bup6okBJdTBbSeXM0nj6HTjliyq+xPho/mTiD52knsJ/+7tFoCz2eZ/WFDIW
J9HoPkeRY0n6NVWYa42oGVdpiCwWcLqunj4i0OV0mrmwyiH9Nh+qwe4Br0qMoSNHV/iZJz6Zcl/I
D40uCkXy8N+Ydb1bxSP9Uo4Yk3HZWg4rJdCrpMx5Hp8xC8esofUN01nnf2Tk0R888KSNys2YEY1T
UB9U8q42dZMRGkjtJCtuUT+z4j7k3vW/8FymVktBkDvR6aW9L7AWY3064RTf2QP1Ta26aw4g3rww
/kfdgib/3pqyRI73OJx8rDydwH7U/9RLDqanq96zVIyfuRs5VhU9ywuSUuaCa5AGAkYJwMn8SHHc
UTmmAZNkyEYEUQPBX/JU0Dur/FawHmwwgnRcY8wI7cwDunc9kx9PJPGRUH7EINiFJASOLRUT/6NP
ZXXHUWy0467FUvYLyA8qlcGwftlde1Tpcf4FXDR9aK8OaWFW9C2AgV/kllCj3KqQkrnfugGzIFfz
DrbDN4OL5UJtOVeQviF65h/YrddgbTI20p5VX4HAwnYpardPg5XLq38NZk7QAe9gVtrWiJkTT7t0
bS6PFvN61o4IeQd2ukJhBM7o25sxGMJLLoIfNGYQlWJf4/Qt0DwKrlQyS8/q/NSWJx1KImcaGlUC
Vq9mluSbxO67nrFx64Ds6fvIsArdisxNiTrBpW9WmAaSljNT2K9snQL0fLtCfyJgbnoyNeMhNXKU
pwoNPfZ+yOMX3p5W0nTtzZaJ3NxmC6mG0Q36gsAych+j1hTwvVmyXloNAr9i/wgsD4BgPaulLJD8
Kn+eUvpEUPaUw17Iz428kD1HK867So82Tu+nMW/LqIn48b2YDIwAPzFGevxL4nnNkfG8C5PdxJ5U
wxH+jfuXByAoGWLsLc7S8JjKZgaQS2LZ5Wc+W1IkhTY90c1kkoavh5+jFM9rsZxN1i9UADRnntlV
fG4RtUQ13ij7ThpmieR3fx/evGjFduD871A3HReYIo/8/CHejAE731q1GY6MLwnnqjrpZ6qtwi5s
Ex8RPN79TJRX0zY5u+sCbxyV7ih5ap09KS11C9KJpkQM/c6KUzA5RtIImbWtybe/mUSKyQlBC+eH
hTdTf9vie3XscNSTq3BpAbDcMYgvtFjHpAOq8qVPzumdp55zmvwYXzong8O8+GaRKBawOwqhExya
sTfzeIeRO9Pa6gKD6RqDW4hjx2fdS0I11fTqd93gRW+EJo2AMgE/moBVStu4cPefvnS2PsCDXOXg
/6b5INHzGEfypSgUa7b9sla/N3I7EMfH2qzoD64yF5Z4+bZW63fgSpnEGk1fiErNYs5vgnNVcCBL
uX+ZYVge6zPKCOggkuGiGEoOOcwr8K8hDGH8utdToJouGc2LtuB1LDMR5unptz6c66YVRnL5Wm/a
i5OjgMYyHHzoUiV+UTJZPvjeEukfizSYpiw9kiiedAvQWDyoYcBndr2nWYWTa+kO55/UvgBEBV4A
gB5VmKH3tyBFeOnE+cdpH/dColSUs0GlZPbzMEV8/O+wCOaTJNpvTZHcBlqN4z6mX6h1NKJwA774
RE7f9RrqoiLH00zmxw3Fjsk9AF00Eb8Y2IB0QWza6ekBfuM/aj7JCgO2hb0OSRpOWwJZs6ykVzN3
KJCtwnaOgmJXUw6CZUspzgDGVKg3vZmdk8xUtpPAnI8XiRhMQ8vsJHPlvOXL0uyP2be4hFL+3K4/
+mm9wvbiRgfGg26HY0nljeaU5hvWjkKbl8d0go3jFDBLh+il+mPdKnsu4og9f7GE1ZPyfnRUeSOg
8Db1je3kynCdjjzFIctCjjGj2mz2G52GnDqhV+9bAgssAhoI3rHSaWVt9eS4jgkxRaG7Z7KIjEss
tHAw2EGZ8fel/zTVcZ5SPSMkceGhFG1xGM535zzcspAFrUdYTrcytP/zcUWrMSa+t+Vgi7BfH96P
2GXuZrLdq7L8TS0KVHvplq1Y+hyn+LFGttidbKWulqWl+aRJvzlXtn780gKZoQESsSatuHOFth/W
UO4CUcfkOnHlQnYmG+RtxCNJ/CLk+At/0hhoOH9kIbGJhjPkKqSBu9/4SwKmKR3g0KcLWuxBBHkG
1D6HSx7hrniXYNqJAidfUmAEeWJYu/K0k29YegG5xuydsvs63EuLT3GhDZGV5eR1QlNA1D1LDqOV
irz7GjaUpA8j+0C9Q+FpgIrP8ySicJZaNLWCqd6Kkb3S4zfJ5yYXX/uAwZu6SFdOINjjQUUnBz33
XP+UZNZd2Fwf57xqM2yzSBQNROlproGXakQVO6y73wBCCdVN0RiF7DAjtYlo26rbg2dpWF9Jirpf
0MfQ0qnGuLJ9XcoNsZ8uE2A6K0Hw6L/EmXq1qRuGyNliIYwSXi0BHOo1ixkHw2w9hI/h8nQZ2P7+
WUuf8gtkhE13fGt/AQ3CFfRxXA3ice6RoKktu5lJeRV3JvLBpJm2y9icd5OBO1et36xczcCFTiPx
fz5KFdfaYYgSEznHTkaOi+nVOw+wVXEaaLJqvcpAfk6EDnb1oKHn3DoOfShWaUc93SOCJX/AxXAk
7/hQNrqIp/NlJdtXRj+c8mtOjGVzN3MgJmZ5DUSzeWWZ/iLZ2W5wvJgNn9rp48p+Zt+/dL4Ua4kW
rlf6K4Udt3L9/2l0HHH2MuYeeGCy+14WgkCswgnRI+UiLa1RwmaiAAIJ6tGJALvHPHZY+poov1Wu
GpIFTSF5V20q85eoOAJs/8StMAT8rYHh0+pcSKHzvG5PFiSWXp2hwJpS7FVTyyhX0YYt2w+Gzs0+
1UTbxL26CGNIsKQflor7uE8MulaDMkvoI8No+Y9rNBu46pPdf6a3ry6HfoAmpPfpTi3Trcz/jbjD
moj0B26RB8pvxOdexzq2BmcFm+HlENzlmQ+mtKFSrdJvE3+IiXtiGAbigAg2lJ3MJY7qRihWqLEH
mdSfTWQsiqsGXY5qDJiURjpe48gVtuE684BkDN0e8OZ/VTwqdG3+tPYOwrC72t3q7dNQe0SFxLbi
WdoYjs6/4xYOy8Phhs2G9j8Fj8iVA33vElw9preFWRpcaX1Je6qXTnePInXum+TmCIzRfWGhSXP1
IB8LJIRlZwYs4Sn6uQHg9Qwl7t2U8v4luE3RvkX7owz8H/uRmonlZNvWjsCLBf+qYSfHxtyGm3tm
CmwrQYga3XQw71bYD6SWC6P4HmGxeYPWIhCl3gjDHsezbBgg4LnyTEHcALGoY1GfRkl+dmUvE4+o
9RcMl6Zq0If4b1Gl78lrMkd4lOc9eCW6ZNwyanh4mbSsaFwc8YQOXxxatG6nX8tVAvZZMfeBcccl
1JgkMIyYe7iDbio83nSv+i0aBzNFcenrMyeL9TnAzYgJIYxi0ATF/49khlxYf0+UhayOf9E4e0yt
paWDDnRadxSRsvBaZmIFqf0i7ah7BU0+76lbmCez6NFgf7PSy0yHl4kUAQvQYifYgc+J8rtlaEDR
q4uXAfvgj/PcW1rANfJ0DAT1fB49UEgBZT0fGr8yaADj/4gav4CEtP36iuS+lGE9v7O8L2kfc4Y8
z0ycUi95eSeUJN40LmS7XO5jeTydL0f//gRkEidaBf1f7/YZF4g69OgxnOTu/rmT9ap2sGY7J0PN
PBbt2eHI8BuSuTFCLXSbpNSFIveHNl4QJH98LX8KAo7sthEAClgIXNKkgH6Q7LqKRqFXo0iPctSl
4rY5OY03BHH+FK779nDt2z/RJoXVc/GGGmp9Cf3kc/HOJKNnqAYCqogyHfzTkFAAn5ZOBBCexE0s
SQrmfe0M2UIKru04fIwKfgEvhPcy/yMR99JT323XxNIyx8y3FtpAdLC5Y38JJ2pFxtfl8yrxRln2
AdXxFYy3Hb7Am+M/TK1TOz7RMuzcAj7WUBPV+3DWTxi/xEseqiinMUDd3R1ZD80hizbpvwybiPXM
OzQJqQKF3E/03BUBySuev8MqIZ5PM1AbQLmm7XAs9ZHc113m+mMpiGxWPBeXt4/RPHQ6ZJbapzeD
1pQXRcAGyt4pllrc1ZdlxaGpM5uARdxQmXi1HI7FM2Muwpwaby6GC/p4qEmtAOpJ1WA7HgzXhyA6
2vC6zd/YwGfyFg4jas99bC9sWGHox1elBq1rRESpmoTPXv9XygmxWGrSvhB/B4eE/AaKuJLzgB7u
MP96cmIEEztMe3LQFWsgybcXbd7L00g3OQMNMTXC48Gp8y1P8Dq270dq1f+N7GdB9+6+FyBG0VXh
CbEg+r+K32dS1xv7DYSOBIcwPx4wka1Iuuin545ouhsiuBoeM7WGSuIBd4pVl5y1zYqfHMNhhjMv
zW7TM5MjkOrUdPm8ppS57+g2vBWZuUPtabf/kclubvwiKQtz83CSQ/KDz6X20qCaXdOoXa2CmZOd
1I3ETH9EgWcwEKNLgJldUnSPU6cwh4sqInr72nEXxdmIzxz1p/vU2l3soGdU2pBeIo4Vs5bv9fyi
PdtKw63YO8sa6PQrD4He4vvZJhCb/o22izqXCcbPBGTOKk7Sra+AkqB/9QjbmyPKWQP7DYBpMD2M
V+8URmoZ1w39SlFyXiUi9r2tsqIvetEBUj3XA7QKRbrYjMUzaAfDYu9Q8vYhl2LxmT1CuI50WAoa
S77aQw51/qTXIxdy2dRvtuhbAic737uRqJ+yfcY7yTZwMtdFTSJKu573qyGG5rYm87Rl5gfe7OHu
0ptqsCZismTzGg9VNOGjEERr4qJa84+q/E+VxcCC4AS5GJE/UPvOCw4clKokTtXCnEA00jnURpxV
mKu1P0SMxhejRNeo13F3yNyvo/dkVv02FBVcfc0nvmVF/YhzCVlGZhir5e81EWZEFE71L4prUTFv
NfztPhGyOmvwCHhqrw4UUFCAr/OWWEW6RAli2ARTMJxINTGC0eAifW9Ec/e+rEHMXsMYH9hm9TcS
obhTqjZuA69gmOgKsFEVdjh18LFLxRb5LSTSEQUd55q1Tjolb05xTL/0wtlO3jOR8RwGl2zfaMjg
7UdwGGb1W4RxUfDzzCbSYuYE84I+J/qfWpOgNclO28/I0VKNeXWeSnNj3dMwFNuyjSKgtKX10GBz
MbJ+3RDD35IR0QfKYgaWdBxaCFsiGw5bhkx7Q4An2LY2/qCXAO1TnUaxHvMYeGYWIU4hcIA+p/B7
GxeiL/DQjAertcOyyzAubSxKXTfb6wzs3Iz5AEtiKcFHMrxQc4TDSJ2gQ1KE0fKqVlaS800yUsPx
UhNzGx7wZL+EAn0Y6kLRc7AmnlHlgkC4/3OXmmsqJ1AStVTRfLpQiYPH/enSDpSsBA4kaboTnEDP
KbJed4SxCFRpyZOCW7ejvuRF4PX7tbADBOER3y7Xl6z/JkuaW1sTYG2iy+bhFyLveYXIF5yyVkwD
T4Jm3wUillucRw9fH1vlkywMrIykSmHlX2oGkv3nYmmYJ8awTDWWOJKms8UW1fx1TmRfi33OlNl9
YRRgUNzVwe+dsx8MlPFaIJcLFFbm5yXPCdFLJS3SIwIw6cP7tJNDoZZ1xEX/vL36PHinc5ONOtni
tjOLKRai80k8W9mqo8GyKTv8wMyQYLrD59hOO6Ovb+aqyzUtPw8Qr9XflcrjVOiKgMyscqNdny9A
PplIJskR1bahSweouvA9l/aDrV7SQ8sclBISk1TFGfD68FXF6r78piXntaveLW0EGp9Og7idVAfb
1moh6RB4Z5D6YxY6kQiisoaBErDYwo73D5+9ULixNm6Bvw0nz8oXgf8it/z2FCgbPE/vp3a8FYsp
hXjcKl92NJRy7d0afHBr4sIw6gtCu56IudZwRWKRLAdMtTyQLM3U+KHJAw3nBfFcYUU3c2E/4mqX
9hlU5p4mjahSMaS8RUfLGBEOS+TsX6aFf7uQze/z5pjsNVgDT2MbWlu0yZKzLFCms/0mJ+oluvvD
+HdaA/TmOSv+L3iSiLJRdnxT6xr2jYKlR2LDH0iMUJ++3Gcf3Ms5nHFCPK/gd8JXAfur5HuU6of5
q5UPQvrVkLLnWQ7MSGxOhgDJcF3jhR6e18JyQvtR039pKE9ge1ODy1hmvNYtQQzdxbp4af2WDgO3
5Hg9g8Ya3J/1R/A7Dw82u9HQyFCwBos/rCpVnNrGr2uNczQCpBCjrEO/94sg2U50pOFn+vsRJYVK
hHysc5zhws11Hr3MUGRWYv0ScyFaQE9XAIvTunRKC992Y9pL78u5wCCxmYDUdrENzgC3qpBD4B6i
UbOeg4HJoA5fDs4CkNPC+lsPkkVAMGbfOFs3mn+6BsRqryVJbtuV1dU+CNe5iWC3M8FwBY44S0vg
QoIv0invoxn5sn9bBQoMVybEs8pu+iyPWtI8GTyVkFPPH1hOMW0Nao5UJbFbWYuTPm5anKDyUsne
mIYQcbG9foLuskzt9gITrsWyk1ApoovKQB2L854oXBf8ZCzZQ1EOAN4SSfHVoWFf5cYdxiG+nKHq
47/Wac5YXZFkSf9GGoJSm3APXQPmS+98YXMw6uE7amou5obUuOmknbMdN5ppjOkIMtxDI6fuUVNp
HmzBXuMHMEhOc7+N0RJ9ELDon2S3Rw+96WX3ZpyCLw1wlSzkoT728ty8zFAt4ViKCm+IkN2cJUj6
/HMLqM22FBnaKwRxmC1oKw5qAbXtsQ2i5uCHGCTXjJUUEWtcLmy/4SoZBb6LQDNK7Z2YUh/7SPPb
7NEonkR9DQ8zeVm4rUZQL1qOHnM8PDJXIXegCveYD9J7y4XiKPYN1NhB2QpXkXA4vLnpWrxRNUy5
sEIXT4/6PzWS0z0Ioq0Xx8Ck2njtnu0a2ywcHna1vay7KNucYjUa3keKn+8Q0xO8p7pCQ/F+M1OT
eCgP/KY0WN+XdamnenlhofC4Dn88naB+EsAD7ULEc0R2Y3QCsresCRWGlnRY/SkwZEJcg8Y3KThP
NJrlDg5P/T1LiDybGJvxqcTIFaDsfaNb0MN4/Ljewy5Mk8uI8qeeZ72kNkcMPvvrJIfDS0dOkvvx
dMeStr6MPawZw9E0IYAcHTBZMWzbdxPnAl7WJ31/KkKwsBH9oTjsKd6Po7CiPf4ZYSG28fQbHi0q
yQd3QIpY7wf3/lXU1LJlpRqzEJUZVH+M8vRxrQTkUn3vWZn1zxOQtUaxw1U4zwzyvMOuI8gHRlZz
Q728tpLUzUSecuUXhekH5C4Do9vqsHBQc6QvuEQlKrJW9RW0xy7BzyWCRCdfs9tnfE6NVs6t2KWV
pSKIeflyNBrDyJe1ZaRK4u55+3JR9+3teoUcHkvaoSS8ByLH3yoAo9OOeJRKBF+yGG2ju8PJ2b5W
IVgST8pst5qTWii3DBMm5aE5pCM6xEJsSGhx1pckCSWwxRXLBAQiQmGsBmO7M34GZgyC7xtKcddd
c9Gw1Os52Qysu5qnLAoBxp88M8PwGBd3gOcI+xI/+ee3OEXZSf7mlO7TZvISI4yDHJFc6t5M5i3S
/VqOQ5svPziR7bfKTSkZQWuz0ivFCJ09gRs4hNJgDnizR7/yWmD0gov7rmlRO9/dZPPkCSngPb3K
7JNqdpMVcKad1tGSHoS754SmR6+Yx9Bj1RrcfLlxM0Knr8KlewCQrH5QdHDqF0lDOZrhv0PJFvti
jrnJXEjLoW5YySVNtTQs4UAzQSKFDiHrcplLTx1Xe32aG6tvxgT5rZcKC3O24VERxwQPbw+oHnlO
DxAdfKP8+yKMzbGRODjqv8DKmLpdNsGobXkZtUH1oEXqh0dHbJZKM+Gpyp3/gEnFd1L89Mu9+EnX
uVhFRntX/brIWzd/bouB3g89/XNbg05P4yXch35Tscr+ihMyWknmbVGEEnwUF8y4pLd4WxW93O5A
5cGcbO5NNoEZLhT6jlRhtubKAfvEV6oGSmtd24cej9tttwth38nrE8B8tcALQNpItFtGKz3F9UIp
CBbiybOeNa03IHvzBC2hocZAP2WIP4lwBxG3ZlpZ5/CpPE1gV9Y/0736SlyBAkcgEVc1J/FKxlor
JrvRp5aGRZ6bOEIes/lPAVMf2utYREibYc6MbxIqeiHFczWt8oLPURSK8JAfAqhM0sKiGyMH1Uqs
NBQJ+/9XiB6JIu3/lWmNJCad1mNdQZDAOOFFs/J3XndW0OltLAPpGpQZTLu8Sq3PfpXsqRYPWK5L
Y+V3JsmGnK3pG3Lf9rcx46ZSWDPdTOZbDpAGSbjRKIbKGS7dT0160AsgPRHSQx1qx7UwVJFRE1eT
jHewS2BvfC2NsvaCa1PktMCfZqW8jWEX/fCvHqv1ozqRVPoIB5jW7Qp2bCIHET7fn/eWpc5UY9Vn
yKgyt4mqr1R3ONPe6kGoego/3h4IkXudpKb+Ue9FwRSkHqPx8buzGr8j5T1pGwsYgygAFXUf0ChR
f5YIUi7M3znqZpMDphEFDOoyq6grN/8cx9ICWjS9l3ijwUSTgjftZ8owGGxJYtIRCy+6Suj5Mcpe
Xkr4TOvVDKQJQr6iNXsQo/bzms/e91SFgxZOH4ly6MgVDA1WSSLf4cCcf0j/uNnXKemVcb5lQLds
Y5wz96lBITiVUsUNQIusfsU607I5Hl+dlCNg5d5+Q0NlLpogy6tVUQsoIWGxlDSPI6MzM64lbRLS
43gQ/ugMkTt7coLg8Gn8cxrSciztzFNKXY2uiaCMkuMJ3sXJQyQmiaonOJRKh6qxN+7H2GSsI1uf
9sMyPU9QELxaAm3szcOyuvRZ8lGyFws+Bheh/Yl+ePChaSrno6VjLjrjqKrrDLt6JozbT5Ie/H38
FPtN3CR0pYXwEcC+nDa2E7QqahouOR2G6HkbT4HvhjFgLh0gyLd8zCpQDjjzGGIujEpE9bzQuI6E
Q5ZAHU61XnN1roeHfNhQ19OMYsoA4uDxaqFItjN2e5H0fi6WMm8xDDj6zJdUoy8RK+hu6giOf/oM
PWFGTUkrjQ2gKNd6EXB0rbXy3VNRbNEWODWNLV7wTDJL5zWIIyIUlaPqFPQXXC9v45jxsF3yW0eE
sKQNTV7QgQW0syp3k/5Z0VAXH+Xr6IgsG+E2Yrq0U9hH+noMpi8LDCL06CG0O/pFl9sHJKflLuQd
uh9dhJdkVhpfsARC8Vp5SkFV+OXokoGEO6zyk3rL3vpaAKULCGdscq/LCXtnpX9+ir75BEEsfsID
1JAR/0n2PtHNW3VOgQj7Wvj/Fx9Rdl0plLAYNZURAEsjqQioDD1KWqX/y2n4+uh8bY8n2fF411yF
mHS+1Q6vY6xApngMtSEkr2sSjp+O+Aw+4Yk4b9MQGOONV9VhTRqB2aAG9n1bJTgLjgR+S5bmngKo
CYA+dunOwi+27xJNCm7eLpty/+6zbo8L5/9buOGkx/wCfF03gBK3zVA5kU7op9/nrozHegX0Tgjr
ny4IxJS2m6b8E8XUDb/SaVlsLS4hyPleL8Lp0QpeqZFeSJk3xN0BKOHojimw+1uLWMmakFQH2RNp
QGc5+AV3Kv5QnTUlLW84QXmeeJIrJtAC6nEVV7N9d3MMVQZWYhgw/fesAYqM6xA2ICm8Lnw/gsqs
5VUU/ch8hKEzGMFjb73SKg2BIKn2ZpzNOS5gnddWjJCegNn+XLngvgVXysW3xmHrg0xx7yDf3WoX
pj5TwZ8VsqpyBahFa3vyveAjZKBzhXZmRo1lknRWx03zLz7DjfcfRTE/vD5fcoCTwqp7CYSo/gLE
nIl2WVV66DlfXELkD6OItlWCvnJj6FOzJHAaKFYP/o3wLYnZwPj6+sKgKpJr2Xhpo44UJgM9i0X1
7M6y84kh+mv1erfOf6U2bi0NHVE9pSJDO9uF8WaZ/1FlGh7bROpk9eZiott7/HrHD90WMouNCIqO
Vdv9ODJA0vqQVIrCPbzzCOSmpyYZfT9UiWdy4fukWtI9LHzuulcrCx1ULxUpFtjDBCGAnaGdSMZX
4bsJSZgWvnkoU50sRYC8OoEgcmqqE3HZcbYMsGl1E7cfSs8hfQbyaROD+Ngdy3KohL0/SIu8fsAj
vISYWDXUcgICOq91IlL573+xcUol662fQJRuL3Km2xdawCr4bE6z94KZ4+bNxhL0UobopN3ZO6TD
JUzyPO4kUVivuKyVPauzcmkK9AYPq8mHRvdEZKuIKRyADbPE9yEJHW7HmIRlzmWDCYLS3eQloLgN
PCn1lTSzDAAXrAJBqjlMH72iaPl7F5yveX+GZHn/iG+8q36rSAzEOciGQ7VRKeIsGsECYKN/uE4W
+odvHcJgYaNCZgYkFlMC0HckLhr4DAlNozSrQxfg1R2bxuqJLXMHmIAYMdikdbWWdXewHzmOIJut
cELU6E4DW+ZTYeZ5IFLQxJDRMFrvd3cghrjCFZAOxIY72LjkGmrnX+n/w2WL1/06gTdx7TxXTxFb
HW3MZjD/mOQ4FxtrjmM+7T+lGeyRE579roWHp+y2bW3z4PpRhK/EH5X6B1eMGyqDosfli8Fr0Y+f
QBl7jqY/hyBG6Xu7HkyRt9dxsDrBjYUV+pnbkP0fa6wa6qpII470yaXXe4MG1B9igvjuQSbSLjJg
++SjMlwVd7AIgkz0XujJOC1s3GePhMKjzRYtL9QzdJBV49ygAsr1gx2XjtxD1TvJc4+sdNThFGwh
am+d7hi3h59GL3GUUPs92P8iHPC+HLztdPsKPf1LU4j8APVnngPEHXt1BmaCVqDPt1Zy1oCvzW2b
BTZem9eCgnioytZOgJtKlvtcuCYCbYZ1e2Yvklh2Kcwd3vUekYcxeAYldgrL0vtxKbKZ+4/bmhty
VvhjFPIrUJ91mmnnl0WfgLJz3WGP0Uha6IhXvx+4xH/9KC7DQQg7Z8RBsl7I+jOrXymGXlqFXTAO
/jXCbXL1CFD2IGucAZ+zsfckqB5qnXjbM36jl/56e2jNas+BGdJSjGUkxPXAaWEhANguTFdiSxdf
l22ezRVvniYV3h73oEv1c19WRi42IJVXZcicjvTOvAtWW3ke47SzjhhFSuxwZitgzAUP2xREtReZ
I3CgQrKXW9BMRAjEEUCSDX368GgTWnm0YTYS2zmF4DCTrakD34sWCeMs5wn4fhhpqsev6cY25rt5
jF8FQ7+oiqSxeZTIK6BwPRRobrUNB/IGa9KkJCKmN9RirUhplpfyVxzkEBySBAME7oQVV5tcY3Nr
d71T9jZ3WbJLEHkJas1gxwPdh0sKC3u+4IEzGN6bWqn6cEFFoN5hzHiRSjqyGY6snm5Pz8oO14Zl
Ll5Mpa7E4u30xR+y9GRecrOD+qa/UPbM17aWvAJASaGKkIevqEkh6Jqz5peM/WvSAY4SsAs+9nL4
4dVMbgprj1Rxg2MO9RCd6ofkrXgy/cZnXtsY2nxucy35qLFjmtw/JzYXwXXVDaJ4mq1rfWWUExUL
ZPZ79qlVelNrjFQt8WiozQJhP8ncw/fu20DoW8D52+Nx0pX3A0/uaKNt3JFEqEZyy4XxP8TcX46L
2qZpURUf72t9KajfXyy+wLCD0g1tNJZHPbVmfYFmS9dWXyQyNKvBJVg4VOMpyFqa1LB4xfETdEUI
qM0LCnsbEEnY8Q0kmZKiWnX0tUPbcihXiCBnsYuXNQzm7M6WVnhQ6dwRPEJ9maU19HCatT7hOcE9
jCgPnbsrrIJDLCkvQNx9Px1bHK43p7+fg2yvaX3LKwfqbkCNpPPUJrXe/R0RiSNhmUsCxj3iaK2t
qU98Y0TLR4DDIW7q713j07qlySddgYZ5FoQHZFPpNQWMcFydxxqZ2X/ihnWbdJxsJWx/LU4BXh0F
Ypyh3P9xJytEzfuwuQzOWAwRQwIDB60He1rVyyJXJ1S89jXYOY+4fcF9y/iIWeCptRDfG6RCdmI6
6/M9UFDuxKpkPalSzEBvsP7kKUAmzbRmJX2LPkraJDNrerBTn0y4UFqsvbTZBGR/pS9KRUD278N4
R5lFjQIZPeBODffNSuaQ4kzx4xt1d/cFPTbfUOG9y5Fu3796zey5iUmhQ+TAozhZje28iJR+3bdA
MVEhryK7iOIAq6mYX+GvSYHWfghsL2Gc7gn02Au7k7YzIwuT65vCbk48mrMa3qkasitVDH7DGnQO
7dXPEthrs5d65HVxsEaS3UhSQ4L1R9eI8mO5c/p9HGMxQ0WRJ5Z3QvsZUvJJUIQNyD8gmxKD8gwk
HLTdDEGE2JrJZmjAGvk6g7DOhApas1psAzyTiiYMkF0lyAEJsqVtQXp5xLFAi67rc0TrRMAED+ae
s4rlKCANiqeJfjpIavIw7GhyaRq6LkOwUEAoWXtGUTnBC8lSfev2v/YYH4mruhStjVLyhanEUKeQ
vmj4Xi8gfcZp+QE1bzYckWPmXzXdokmWfUOqNk6aNvEH/y0v5BBc4zpjkZaZYb7ykN1shkE9k4BF
3R/hW7Td1dIyf0IUv7yMl0WW1btE0Kp2PJDRXmEwMEuclX2VKZNpnYcxn4fEf4MMMp13GnR2Z0pD
3ZqTxZKNAF+Iqvg3Tcv5A7H9du33NIqC6d8wKyzuxPV22h4bH4vHj/yNSFOGXQ3StRjrxxltrRwL
M6peSYFzq7qch5sMEEzxmkt563G98ZVwZJ52YQCxA2qOroKSosXLBoyO2gO08YVSArWZAvoZiL0n
Zs7btO8xS20X9Rjjza6nMWOZ4HxKK0o2rEbkFOtK6pw3kwp9Xmn1X7/SOXBF3j/Ow9HvnIwHL876
KPvRWTNN1gQDy5DYR0TDhQSXUjXgk6DBAPQWS3X/her+m2JbrXSeQeSDx3/3HqwmCuBlU1A9xSc8
SfBRscrRxmncam4WcfnCfWDPc6yhO4YMAx0oJCKsgbcndiMylyFvmDl/xHE/Y6SV9XqlStM/BNNk
eJ4qmV4MpU/UM7bd2UdtxJcHnzp+LrjEYWQuZNepwzsYh/epURVyUWCYhfHy6MjwAgDuRUPhtQuA
ZEKkrUUd+S6dfPJvYY8N1M3jaBbajw9oFLp0hUopkDuMPIdIXzqE8T8e/z7i3aQER90IRBtwTHgn
v5njUCod9efvSnLi0YgYZTUWUAbPWlsnHuXDKpXIbrabRaKngH0uWpbTuKXNfkmr6VbhsaeNedTi
pMYrlLnzZThY3TGNzIcSq8btt56lUdgGbxABrWgdfxd1+wcHFjkNYnZH52K8K/2KaAOQG7wPGLyv
Ur05dieAsg/5Ot4s4LkZBjbJn+JnsuGEwOZOL0vaHlEQUSuInnp+vvaUQ/QghJGIIHTJYqEillDS
ugj3m67TcRiJTJS+wdPfFnhEmt6l+gSyGOVuNtPYTvUI6gILNuEv/RGV7WOTvxRpirOtgnSH0WFD
t0kmw+/qMqMvLSyhXXtvXuySmQn+intWPYwwmHc+GG3YpgBP/4WQNNbgJitYaAdYoHvD/NEq1MNZ
qGixlMpoLjNLH2AKRhnzx8I+DgxULVhKrXx/AijrCNyllld0/K4VAys/wGjW0WtWDpNEEZzjUscP
ZnQ8yo2TBFZ6+lZMvzzgznBMJsfzZjo8GoiIcm585GETQLEMx4eQGL8DNGYJHPFKYhAfBzpVV+Mx
/BdlzjDbbIjgeDXmVz9CEC2saZP94d1MIOMOAMTTwIrapVt2WKaZB/OVJKj26l2AE9R+11ibeP65
i99pOpI3viUXAH0Tjs0sd2fNS9KpqqZM/wLzukxvN2fwtzOSA3JPP8MZrtKFOYt8sRc0yFJ2Kp4Z
hf4aazRC9W2vHADwsKK3KjERi52w35K/D/+dE3rb+enhM+6qArmxjRBLuBC5E+jGsVGCI1wQqxyi
jwuvO049dtqpQ0aGlVty/MAuBfCjOUXSGi4nYK17ByNnsCZkRl6Enyhuq7QyqazdPv99AhPcQEOI
9ycoNnaxE+Qi2z2Q/2VeCylPITqrxr2mOdiB1Aucz6RqHmkWZL8Jw0hSn6KM4gfbpMBYNeA6KOQ/
Z06Al6UBsX4ij9Ug5ioe/KoaC3QMiEdEDUJTHbJ7em3GGrS+pHhzTT35VnX+vAIbfJ8WnPGmv3BS
1LUxgcRp5likD/VPnUwKcv8pQnW/8NB98yowadx2Y7fqXp9XaNpgpOvGyf/zw1TAU4V5l5n+xWVr
Va+FzKkVxCdPdNjrkNLmrC8nKLg6QHjs10UiJhItAQNO6cYYMGFLWTmfq9DtJBDjw5LBGlREYK+I
Zy3KgGidC+CtFYm8UlTXQxkax5wqwRWqg0zeau7gdEJookOEm5ngksnxZuI0q04/m30uJL5dbEI5
LTLhTncmaNzrSIvS2YJvjEX/lJnh/h+Q8r9n2dIi/qpHUNARFm+NoVwApzOo0i109pdkRhfzpS/u
NxfAPu5HaZPnPFfKP0oXECtO0Q4GOQppgC5yQu+RuvBQODbcPH+XD/6MSnh00itFJUzebu3HlyHs
+Ifj7ezLeVvZxn5r1cgpFa4RE4NZkxgIxS7j3MyKYOSGcK69WZ8qOSfyvCBPA+QugNNI7FWhIU4D
XMCjRlodctUwi1QqIXTbA+w8fRehPSn20vpx+eT0iUF6Vp3KgTbyVQITFH0BsmK3RKOxgT7/Yc3t
UdjoHf74gcP84BDfMMcZRNBBog0zcWJ494TZLF+DdDkOBlPkownXEiwaC3KF0uneBhFvt+2Yzg7A
Uam5y61Felmx7kEGZjGnvUamT8rcz8crwUX6qNZZ1FD+eNtNLynu+RfPZd7xCAFtXVZfZt/6wjtC
7vuUe+WNbdIYJ/NTRzTc6NlTw7ZMaM1WHacExKbJlOzVNIkCzV8oQhUgUb0NrgMxcBL3gA+HGKrY
bhXbJ99MSqdXo9D6yLCH2DgWqqfd1QaQewSkSdrxlfJgkjYZKRys6YTVLbALGNyAV6fYayYXe9ll
5pArDxOXdhKA7MR0M7O+DjprmWjhostnSk8+MCJ1U1DgKb1ZdVJOCK7Ge2A9Ms4mxTM8QKy7c/rF
VCwHiqw1hd+05IqkbcBOb3JwssoeB+NeqACQYjAJ0gwpZSGnCE/j5tEkK3RZGsS8VYkeHvvzn1BX
O6gjG6C3AjRdE61nWxpnicB6w8hFIaY0QCAd9JZq1GGlpjlUiNl8s/f/FGUpCpU6/rOvdht1P3Kp
TAoBnu7kopLpFQWd+49G8+UZ0N+yhOScWaAEEzasewcS5qPR1kC9OfVPoNi0e3Ykdr95Sgxx/1Kk
HRTls1jLYDeEBUFGf1HDa1ts7hMJXhiFkoEt6XyfGgk89NsM+gGCQIyoP3Az/ycHwjhLHYkOejJB
hhkLSlzIGzRSB/2RzYcOuj1bMQLn666z9aEYcI/CvS9I9xs37/DMVo5LA3NREHWCzhnBDBnDUBQY
F0EqoqorUKZI/dG8Ec6UfhszQ8WHlJC6K8O2usv3mqE9NpyxeRgIYZA7Wa3OkVr3Skg0EBQ6Rqhy
XMqt4X6UMQewuR9xf+BQHdQlH8G2j81CKAjuEsjqib2AcZCa0OujNu05wBJTx6KnN+q9ecvCqaPB
UKTii31EECDPAslI5FrQmHAeSwfe8+PNJXPpT6V93C/aoyZz4EytctipKgwZK0YlcW3QAHhP5sSd
9+eQVC2PtHAiYjZUWgfTTUtWn7ua9LQrENtNhUQ28UbAWea1QlPhOXzXpEdEtdgtn0bwPG6JDW0V
YXgjE+h1OWniXx5P2Fj0KNuej/lPrP6TF/vppYu3g/5zidLf0jq0hDT+c4vk4t9EDMn0IKi+2eoe
RZEWzUILldmz2zuHKEnrK26frlNf64eFIowduOMLaKCgV0D2fuSEQbfDkqKLZCTn1XKmG2svP9ov
NTgCsiUes8JZ4LKkgzgsHENLJEOWoJZ54ECIJbylXfSHCwnw+V3+CiCzoZxAL/VSoKQnPS2/iyuQ
M5WtpSONHhEhZ6QSk7SVJjnSS6ZJjk7AdfohxQQmkhTiMDglJvuWmaH8Q6IDlT6O/jN4cqhTrNSj
J9W/YpWwD47SmubhsJs032UDcqU1Fv0qJY1I7tMFcHJGP9xifw6eFrQRftGNm8jrhUjAZLJCowdN
Q+P+4+DCIoxUYmx1vaf83SosQ4xubhtuf/uVJIlH6lO7eTnyF9C5uv3NkgxMn4SI4ijeC7BLuXgJ
9nD50iCMcNoCmWYnNCMeUZBlQ8+hK5fXz75jlZ7i7eXmvuKiyAsCw7hrGQSXo4YjNH4eenRspbLV
Oa9HrbK5SA5uQVkvyt1r4J8wL5AyX0u/sc87u82wQVtfY21sw6fhrcSEotAa6fHGJYTQkMzgNWVa
JLHLvUe3TkyYRjr4FK5qBuLigclpHSheZAi/xCWLfJSUdEvyA7PWGLC8f0LUIZ5wBn0EPOEhReR/
1H7/MRiU0Qt+CvqgCNoWyC975lc39PjVnRDj5TH+4LHjHd/LiTQNSOxMYR54QjOzko9PYNqT6Try
zJv8sgWm4ip0Wgebx5hCK/Jt/8kqjV9L2JxT97Cr/q2IbIKaLRWTUec9hYq9NHeXn/Nnve42Zviq
ES8sBw0LCPPs5vFh+PaqFuCv5A/CtGeIQKFSc+n+zfZTIDYwiDcFYdDPAgGT3pjI/ZJuhaIHgsOI
uyHBNhssiz99GbRkZ7teR0bsK6KwQiAxYbCr6fZj2/PcKQ1UM7Q9JbneGStNi/XIsoppboxssf5w
gr5PEj2dirpNu0vveCWPgdQqt7vUAEec59AIXZQipM5T7sEtuB+VGjKmp8sertX2V9nkV6zxkp2r
dsoMdWVoO2EAIJS9YLZX0TibBk4QLlzrUX644+OLNcKJjHaCpPaEoWfE4F0riEo+E3gafpo6FqHf
6bRG9yU57F+j4Ws5IHZttGOON1NsNrjf9Rwo7fyRqZ3wJKIW8NqbNw6NfqpgrRtYsVYzH+PWlQuK
wOI8H4kVlJ5ZVC7lOtFFDGDU1vCjfqcxk9zgxj1u15M3A9IXM7ndCSvMHkQX0CwOjnrVTO0Qkmhc
f0Rq3uFl1pd3stGDEpRVkSw90f/EClPSfHo+bE6aWezW9duqFpTGmuzEjZ6DnyBvu2KSoccXh58y
zm32Hyy964gWIu2oKU49s+ByrZ7RGTKbJmRxKlaFcfU9gm9kOqZuIT1fK1FoeUC7Q2uGI0ugd6NZ
NMhaqKhaPFdLppy1YiXkCwC+mE583NQJnTHpS3HYS00VDSBZ94gwuFG4fJ6n1yHSzxjbPtPdMlbC
T41Lscn29iBYwiVCnFQ9QIyAybW/siqWfsdJqH6yeBXeMxY+p7i6wsg2n8n+hvXzFKvi+x63clAX
tvixnHDPVPDZhvIR7/ElqU4CZp3okZlcUAB4OCnuRCHkfR4hCIlTctu9QBql5BAjcFwmwPrVuMOM
8W0DwKe3goXefSzNvDJOKsRcA0EzitTdfuXBWMheSGmvGm4NpMjbE2KqRpbiC2ri4IL+FGf86qnN
05BOkkB16y543UwKeloO2HS1N3iluYb6BAw7o1sb04IkL40KC2zLSdllu326TNQAmAoFsy6rpvgf
wG/BHicsGjPKsALy9upyhOyov7W3uA+zwvaqy4M6EPJpnfSMbOoA8Bo5z7DCb/hipwg+37r4cC+O
qNjSQxefx8NakZkE+GjoZa+slMCnI7GVJrb8m1NevA8Em5fus1Um0DBRMCojUeqmYjiYc5qNi7aV
rhsQ7NH8Ax2T3VWU+DjdOUNg9W+/e0B5QuSvRS4XP1PjJQiq8Cv+5FKnBgaolcHg4vY9E1HmhG2K
jkq7jHnwI8eAoLvJg1AJQwlaci7FuwMDwjv00LeW9QS7hfS/n49wWObZr8gZBf3jmQ6R7v085jQT
EfAOo6keUghZ9yhnZzavS/lSEC6n8RcURAqpdMxro2iKx0om8ioe4EURKzX0lt5rzOHrygCEccm4
GMOZpysTuk1buAFYr1DPpboadu0wSB9XSoFklYM8riKW36uIxkYAHvdPgR8PFwAfFGs2UfhCmc/o
yKBBXDs5PVW3Q4vuViaWHqDZ1YQI/jiL4op6o0qL4/GCaVCSc88KAuMkxxfujwA5nIqE/elim+LB
hJQInLaLhKXr1OLPy7f4rswIHXJTFqrybLZW/x6RSZys1chyZxDscWLlRoytNB/Z5z4Mi46A5QV4
ExhyHfjD8YMgzY9nB8150MkO9s2PG39yRsunyJlDqPsdSOqruizaRyQAEkyPdjK86LJyLDCbl6u2
ZEAIUzJF5Ec3UebXpXVJJQ8lc0jG2U0D2r0LMtMEEI2w5mXQoZSbR8Qnd2oBcQp250OAxqB2mJ/G
qcqEna1WnAw7r/7u01fLzIqkEMzXyWzBY0w0ZeGkGN06A18b4RsP/sXo/2iNmNgDE52YJWZIU97Z
AEn6/jd7WVViIU9aTCpZ61oU5yRWJhWl/T769Pt17hvf+o6GcgVwsQ5MNwRV0fEe3zB7Eu7RGIeF
buHEsPHtEhjeeXeveEbanh9PrPIG1MwTrSTKO6NlG4gXx4PeLwA31raTbfFIhWGMN/NAzgJx73Wm
Qgp3o33oU6+/tninMfuU+zdM0dask05SWYcM0/+f7tZVWKf3pszXTuD/jSEPBLzHjAYyxXuhjveQ
bgBBJ78ncdK0rVjmHXuJUL++M4e+WT9tQfI+yu/hZZjZUAbP5yk/IDGquRx6fv/rb3AEHLLdJFsb
j81dcqoEYEv8eP8/MVeWrnqtB5/IIAfiXUUCR25nSzUWNR7eREWpVyuJbVwjO6OW5z7niTqDdgnM
A4v+p7Jj9sNNqu0aJHpvkZ0zZ9X7n+n7dbHeJDWlh8Uf/jJBYxWQemyvfdAfmrZ0zS8TEwafPb9o
phWKsT+Q6uUtuxjmDLEncqKXBIedEEuyRYmjqmdk66YSOIKQD7knT5ELTUhkmj+PIvXQxlFnEnfY
ho3f2kfnWifPm4XJ63s4CaKazfHzXJj/TmAZ6PaGg88sXiXAeDNEh/d2YoXzjZMeAbn5e9u2xOzy
Nfu3xRzyG530Esct5lQ3c1VzmrODUXhfncJLkNzrwK9/MS/nV+vbymAuqeTZxine3qxtfb2KoPlk
UUkE/D2RCw4bmjvj2oo7Pku2wXKOnR+3DN5jDjPGtC7gQxGOnWEopN3nUIUO8A263PPSCHxYe4tP
VczM4X+anNBb4RSuE+6+ajwBHyBI1gbXVtjz3/AJLAw7PQ/jdd3wTOC0bYVgkyG+8DVp2Fy/rBAw
gMRSBuvXG0e2+K/vX5VQd3Aitp38LmdV2CVQVAgsps+16fCnT6iDWK2bwHEZLfLMIRum/nOt7Ldj
HpbnPBq/KngUf4vB5jC/MY49ey0z5KI1wrnNTxp0KIiDyDx3FMXsHHyz1zh5MamZQH00JBFT4AA6
Zuh5O+uUhiTGzrPAYBRA758XFg/tREBqETvg9qepdJ1MdSclb25ts15pcADrILACAN6LjCG+W1x0
+2aV4Z0oHRViWrrhfKiKylTDMIlKNiL4Hf6HQqCJpCepyPFysNBRYBYkIzray8zcPaN2dliWZ0qX
mBGc60OE397j6k5sQXLVUiBmxoZidpm8RqNFhM0TpfeWHmXeQcIYneRRzgxe+A6QTD5Dy27luwYD
aYgZjoW64Y52vrfmCrUbJuClJgAt+cmWySAaEQyRKQnPsXqUybTJidrIIxR3EuhoUyDqZTaP9mTo
D3qPfGV84d4MS5lPxQo3kPISxywQvzzMAGaOCUdjdZ6cw4kI2Ur3QEKHh3IjCA2J68D1ACw615PA
3VDYSVhUbL54i0pKRFinyTnNTbtY7w61aFunlRcOYCnIYfL5sg5RD4dLulAkmTISqaJ9swp53TKN
10LP04pjT2aapsM47OmmMWfrtYW7xS1LBHGvY/kAciZWgmCMXBKOkZlLW0HeBAWNlcncI/cHq3xq
/spfIg5bR6iDeVWYxNphI5c8O076pJUvGF2wYO9y147G+Aigf6e9fg4/6ZOpIl+/jnmsURe22NPW
AS3wpTSpgNqvI7e7bAtGgDz5y3782ZEP23f8EZ7tZ8IRGHPLMGL5lRfTquDivFEW5RPIjtg9ifEG
JQP/Vbvt6ymRId/Oo6frq2Fb8Jt26SlLo8GEbefDymYOe3iV26MSvFr816EivExet8f8/BOps90F
ZjBpKQWedBArl5OXLQNDSZuPPfCHiUM5fzDKNW9YNsI3YzLq+cVZaZS52D3WMpp0dszNhxNObyzz
O+VCZvmHR3xY9uyL8fN+Po67IYYtzAKXApao4SIkxXIA/TtHSxdKXyjPzAIa7QNTP3TMetn9JDbW
YKtsZEG0MADPabRdqI6Wxc9pgWZcikh13r3xz/KCS6RryWPPfC8/+48ZSu/M4l8z5+H0TcwVHJwH
4r4H6cLN3LIp0SIrN823zKLTEV6KkVSYDH6LuwuHYfMg2T/A9YC10+NhHi38yo3I5/s2ij2BsZig
PeBa3CKQeg+FFmc6nKULTJjex0m/fJzqnsCh3PpkZTt4tO2jQCbJeG5KWuZrSxMlT/UXJfQXwauo
NGFz1zRXjHt0fnXHgl5Pfec3U0CvDhbhkI+0OB7+0+YrJJ14eWRD58OUmsvss4l+GbkLA86BYHfJ
NqdIX0joagrHgoNr+Re9Vy9sl+eq5la5yUUnXjkC+OiwxExrnrqXfa7FiPzqmv8F5g392PS6FW+d
+VygUAenFRCdzw282fHl+aClrXA/fT8RaKHRWeLVlDFvtelTGNW7VN7iEyfFp8Jg5CPn6QcJBEYb
hpSS6ElG+yJeSriIDnBN6w58RQMM4gqfkMu+T3eoPoWzS3gVW1ysWUdzOkDq/g+1IuAdejx+k3uQ
AdrYJCjZBvk66Yyemk6a5zPTfRDUowSKY048i5FPVTWpZMJip0cO4l2oajpL6ncagnu5g12XKGVk
xhExNkGTaCLwQ61YFfYPo3gU0CUEoKNb4Fcoc05NcOJHrt4k9AUJZ14QCK2fzuiexd022WFdCcU7
YgHLSZG5gWVq2Gh5goimC7lo4M0/J9fjncPplLWpO8LnXfjSwoNI78KR/C7AN4pBJ3telyaK7iwa
LMsDBJ8Ff6/vWckGs7kIU1wialmCecG+Fagfc/WlFK/RZUibF++t0ekHA2Qh2MRJaPvUMAOQLWgT
OHzKckvVY440BzJEov6RSoUNUfHaoyOQrnOPDr+ykgqeDCSIRNUQcG1gYfkDCBrdl1ovj5BNa4or
zm1M4CR/CB76Ii63RdASGxVC4MILMozvohkYYP128LT5O8NXOy+RhTtIzXVwUA5+EGfHMfefhyKC
+HjS0MNrCKzz52es2AVRAeICQmtNuHzQduYqBCSN7KiTfGUII1+6Lst9snmP6hV039VUxXGVqaKh
aLozcWdNpFUlKYIdx/eP3lacwrtnIidw8uO/wkc1//BIGxcq9l/wncrFfq6P9Oqogp8qwK4mNnmu
HxkCGYfj0vB7e2eIzDuBwo19JXb9yEGi16WBzwL1+F5hAIXfoukXntBIyxU/OrRyqLRNsADX63ax
mTyWaidMbCoIKcJjc7WOFdYYSU1EuJ/Kb6V0PphSVOeBLk3tkUHy7qLsl2xt3sRI0Co6docKvWbt
s7fOW7UZrMcqdtMHIbxpF0NiERdmLnxk8gx7ZlW/Pq7EO7amjwwHb1XY2gS260rm3i4USVQEa5dM
25Pf9OVZERYlYdEhyazz9QpOdbjIiFCS3N3uH4+hJtAZTsZZqgkZLyuXqzD4oQPTk8mocEtvg80/
xT6EgiFqtALkz0vjPxa5VRq9L4q8ezj4Jew5EaiZhnXmlI48o+Qz2GeNWFoM0odiCh1yC0tlzX8P
KMdOFSBULtEi8rZC8YvzyTJy+xvoN0cCM4XhjgHuUVGV0vzIF6TGEr3r6XmKfg/RBH0qjZV2bpxP
MkAZnY+1m6wsEvUwt089DXdmu5WHFf6NFvJx4EiAKn4fRicWd6l/Jzy+nzusESQunbfpom5DH+rT
1hebhhdJhXPJYC8l2dBzehijCzEE3ys5HNV2y16NG66Xs72FChyw//C0H+Slj2MrQe9kSkWaLUX4
GRNB0OJFX7jxddW99QQCTDzt0c0egqOknCveAVDEwR7aqT5M2cQ51XiE7kcn1x9YguFDP94y1Lpa
oLhSkuaJD1b+3oZetv0xj4S6mrhJ50vUc/Ywdiav7fLggQo61JHHT0Cl/z3THXyEoWT2togQ6wcS
lMPX2A07bbi9QzxlJ8AoO/W+2awhzZVG6CHQWD1ZAbrIumbOIXJ7L1MDvGyS70Ky7iql99Su4QrT
nNu00JOxts8xpZDQEBidu3iiJ5mkOSBdeF1A+djULIWt0nwYeZxKBd+AQsz/+iFhUU0R4gpIc3qw
FDFvHbGpaO9qE1DA8UkKgS1YjjcU9L33Ljn0ekClH/ydjdRDZFI9DVbpdSX+y9SCqX1cfZKfpCdm
mGMJzDlYte5Y2Vgfvg7MWFY5XycIsDa2ULRorBNXVLt2yaQ4HxbB0UIA9sYFFTaxbnHWSv48hPJt
ESKdTRbK6YOFvfPuEBerP+SgkgCwvAhaJd1c5ylTiPivlhrRkVdS6KdQmP68mb1g4ynSlDmpsgkk
RhzEEbRjMbA7n8/eXXGWiq8LhrX8NNe1Ez7c4CePZOFKlFQtx0M2Oq3RnUulj5/WY/cRcFCrYatb
nGDrmU8scjCtSAkPOJLEhhhxEl506SjQvP7XPRwzxekCnr7d39DhCRIAuxBnXV3XQ7k2sAcpeJ4m
lUwuyn0Nbt19iQIGUUd0vXcGDXb+RzAGE9Mzsd3XDezG7/GtU48VTkZ7x+jkDksJgmGWUsZMa6Ln
VvAMpoMaDmiztEnZ7tEkdDFEkuRkF7uPc1L+Q0VasvAjaZ/AbWYb+whNkfezrXpgmzFM0ExuUZ6M
wBzYzvvw50qrLPoV1zW3fpXVkZfO4D7Vi9NflDQ5EOgLABzWNk083ZvXDV6WCSetB+sjp3+ZGzgo
dLJxJ5HIzIPXA/JVtWOHWVhZHgvCl1smVgEXxdI+eC3lCohDdf3D1N8yeA8JxpEkNP9D6by7XAd+
9QN+hzmNx0DQJLhNgCcmGC5I0ZZwisLgi+tctbNoxfJAjkuKqgoUToEO1f4jgmU4Sh1lebWyZvER
jchQPcUu2QS5sfiiLISdr2OV67SDG/OuW+Rl50Aqkrxgx3WcfMZM69tLhxHKw5eZDRCnW8hL6AZJ
MNRHh6TuqN8dWtiirx8UTgyRR0UjQjpbE0x84KRXa0sRGBUcv9VWRdf6yUEjl7o+UvUxCeo1QAVs
2SXF1hJiRtwbuIgKc5P2h8wJ6SxBga+DawkUVWNZo9KmAWpeeLfryozN6qe0iZFtPUXltA6vbVYd
2BVYbCJigWwTc0h3DZbBK3syY9dP8NhrKG5RDIYiu4dgH4xYT4CftSFolXRq0vURxvyKBdXIDSf3
K966utnjV5IxCtCbYawu/vVFRwSfNWEDTxwV5nbyJxNDyHSUYuL6RaoQcsbb+8P1EypIFYVDzjH7
UgrsoGxElM//XHDIarcptLrUokHCYobGWdl7zzqoSBUWoOQf2MdTPl5F4qw709xIZkG9EHK7CuKu
jcp60xctoK+TnkWl5dOKPYVkUxYCHV9n2UhLKGJldLLczbHW/NA17Ok8x574q1N1qRYMiy9U+IoA
2QBmew4yKVXdU55lVlroPZ9YIsYugQwplmLihmlm5hHkKXjsH64TgIluZ/fFIxWlDVlyFGFVkR0R
TuISH0l4UaDob0S6uZWVOyFDy8bHaDwV6QOHhoOJ3BR937zcnjO7daXcJgRczYsSyndzo00mp+k/
T6dfIkZpt0zYV0OvQOrDuFUts85cizuIl1YQu78eqy79vOV/TQodbXWuiQbBvhVLO7Z1Wf//P37D
Zrjszfl1plALnBSaJQux2zLJHLh6hd2HveJIiuGVbDjg5juL1uGB8ku/0pfEAyMK/Avq28holYTK
AJe9e1zp2DZpUewaiuSESa9VHLAfy/EfUCvb5bRCVQaW3pJ9SY6KTWVI6L5SBStLqiY+gTBTH4tD
4EhsSK4fa3AbTg04N84eBNHIzAFcC8cY8Y/rxolGzKPjadugXNkoIItD0SVKIQBoPkadzSiDCfS0
wDG91iLDk2CzdqXb1PtXKzss41DsvtDwFLVdk+STPRizmwLwTOq9gDNNIXGW49RMEotL0HBUvFMf
oCXFG2+51dTa9KIKO/OrjV4KfkZgxLAofm3JmNVxtqmBurQo7c9Xq4SQZGqoSitFN0z41K1/XME1
bPk12Ix2QReESoushPY5wl1v5nZKGpq0VP4uAxqhUQamqDOHtpdscaAGjDjgej7aVdgz28y740tU
MjZ2Sqx/0tcpDWERonVAEjd8DuGK4d/4wJwG0l+r5PX7AjjeHcQOLoCrYEM5/wv5LqWNGEiySuz7
t+otd8s35cUHXGKV3NY/IEBJx20JtTXQCCV5iFfeFh3f2Q3nihCVDMh7JgeXpg1J6dBPiwtSVvHq
QPhWTYq6Nn+zQikoqXhX0TLG3caTRXRNVVWry6kEnAoe4Sj/wkSfHM+B443y6e2Zw/hUb7APcqOL
zyw56P9LliyZvRzfCD6zvpiIMzNAGoLW9QooUsydbi7dG9IViRL1QLw8XUvRpZVYwYxtIE05arn8
eVhfMwU+/d4j9wNEjNQi08qbCdEWtcKQASzCElAw2zT7vL8OsQKkHYXzFx0z22HuGz6fVzV880IP
FdvcDlC9MlOSTuC+uTFinjQlpu6wMp+WWQnv2sBMmIFjzqWwfqd97252jBynWnsyVVIMF4157y95
ScWJ0tc0gKB3yvlRPWloP+gs2f6REcSGaIlMmMm0Zf0l7t5sKBJgTlwByvVbGjxcEh6Bk8FVEATV
5dHp6DM8qljDRtchq3Zz1CPR4kGA3j3wta1ebjumei0u5abNs+Gas3kt6yvdNo7hLXNayi+gkhUp
X3p72CIfJUvSIv/WspuX6/6OrKuwW5YVNNJtr2g3//LaFJjJg4H/+ZM4DbgpzTRbENbyqalBDcu+
CsLmsYLj6u0iTCNvTQPiuxl/WfA+52jOhWbFKR1Dninou7YrXXTUHvHsm8f8j38QrXplpCDOW6j4
/oSB/5J4BxPh7BfM35iKXSbo65PMNeJbjEIWvUanuqzB4zI3tgX/F+KufJQYgdlC2zeBO5n7/cXc
j3mlVPrkzvJ/wO/Q2EhW9pwBKfnU5EMNevtY5WzW9QFVRxThBr940wsh1LhmFOQvizJNyf11sDIS
KVt5vTY06vzuL3kpH/nKApOHg3yr7eR8/QNcEUgCVpHTI/K3vNiUaA6mFZz65epRE0sG2aO/jEta
FuIqcoIoqW6NrU37sdaA6XGOSK7UpbofH1gXG8rbJ7IXmvBFvV6a6NQU7d8RyksbrW3FqoAhGX+z
MX9DVWh4ll+7kf0vBX3QWI9sgolod2rD4qa9ta3NprJt5XDTKWAK2dsl7wYBATVQ3lOWuxnVcuwe
1Ts3wTTKU43Ab63bxTlUszszb3f0Gfb0TmP5WuqLm/CqkfjvYO7ABxmGFmn/AtzOO+QkfirBWXGn
4lHN3fIfefVKUHqqNdkFOR/An2/+o9qbV1siv/jDKkcFyv0TsrxcTUcvSV5L1jXyZaIbd4rXU1w0
h5CXDfFvjRrCuYPfzsyhtmZaMaoaWkee5H2B/la6few1fOEXL//xIGPJPLrSwmaagfIWB90oDLJ5
XhqKntWr4Hh3DyXMQ8cIHHXN4X5BXFfYW3iiVnGEVI5doXKAi45PW+62PKvynIYADDDtIg0KDbzf
Fo+wy0Hq6Mv8A2/4K5FE7rO3HLgcUmlQxqjLbRE4EwLC43ObR49AaZc5opalmJ2KpJj8lCHW9gk4
CLikUmrRY9LNGvpLyx+iyakW8py5su/Sv060RRLAIAWwr/cSAK4Or1kfv3Q9VQlbchWfEGNUoIDA
i/QO5M40+J7wMV5illQ4sxPzCe/Uy46ucMago7Dfocw5As3MhHSHKcrECXXtTrh1k1ZxNVF6BD7P
U7uJ5DRg+Wi+f4C0XEu/0NzTJgF7CXjKpE0b+qK2dsijJvj/if1IKBJBC2nQP/oHIgTFPlC3hwu9
jbSJyj0Kyn6Gr4ipRlyX900aREkPSv/uoZzGCpyVyIHzZqtAj0n8eIUIXVC6pDfYZsa1RSkPthMs
9gPzR+jyIpXyDYjbPIJQ2ooaWEPWD7M7gH7UZm6b/uEFHMFNMDOZTyVcsazzUDCyRmCoS4oCIobg
oe0iLZJPlBWCQRYDylRcYVR8ETWgW0Ct2vviZ9CugG6Whi0iiwzAflqwXaYVY1Pg9k3tpwIIatPx
ngRgOuQqkFLj8/6V3+irqFKwCSb6rlk1KlehBzv6yosRfWWDmca18JFUhLHR5oZwjTX/9IZpLzWN
Ad2R2l/MoetDsSHp3Ce4FFTlfYH/morh0LUumBDTkhOs8d/dCI6yWWlVyrEj/FP6Q4ZH5T98KJNR
59ItBqtC/YMjBWP65jqbU/PHxB89H8anU+bF2kruLibkK+B5HetGQrXu8SFFmdpkfW6lLZygufui
LPwxfQeoyVNWciulzEIaKQKJ6ySp4O4EJQTgt2Fj1mYg1rdytWDOXePyHUTSCy0Iwom4huJRroVk
8ArxXcPDtRz39yqaJV62d0OAT54TPrA/D9T4HPcU4tVGaWlhP8PcdiZdaXNJSGwIOn4iCCSRFanx
RgfCWV+JzdlAIgx4iaZ+teFYZA/37wQ+VG7VykSJhoyhximuungtlWZrSwE9uz2dKtB1hmGC8uvO
JPyrePQOulOrwHFTHwQbO0StSVSfLsCf6R/cF6Tsm6fKtH2IMc3gdyLN6gqR/zrVSeeMaWjXJy6Z
Bq4UYu9MiCs9VCQAnbXt2C9GxG726BTKb4WjOnr5HRiRL4jh4pxNdYLgwcc22M6rtbZJ9r1kdPNf
AZEOIFoMK2vSy85a4lN6JfBAcT+P9O2N5+HqBVbCIcsakBy9cjND+yo1SwO6fPtHdEF7IgMVedq9
ogLr6Cv1kfLbiZbt8iRMn4jn3fLz1FPtwB28Yi7c6uy/eE75nOyg0EZo3Nye/n07DqKq6+jhmIX6
cdCaIVW12ViIxtHK5tQ4S4X1vYi9l6/klFfCHLbrH7ZmFGVQK2QOBnk4+sdb+Rfx5PjnbrysgEv0
C62xU0cvj35viktydvYTOL04+WLC6pytT5yJ0Mnqb6WbaZdY/2WHpp2H1K5nCHHk0ThZu0g8cNLH
qJs4sAlkYR+H0bo2GQLgT/IB7/OpkkVOPUrMzv9iUd+aFMVrcHNjcAH5yz09D6ON2pQTo0835Ucn
NMN6kMLhv1VOt+jLsqUn6Ege+3awYFaEijRK5S6jgGzai7ufuKIVTkcI08rbt9j4TohJ3Cgcmrqf
3MjHgEIzRd46bb/uzJOH7/HUi1Km89PH/huPNZvYUVebYWB0Cn4NBcKv9r32aIKWmiO7H5ixAewi
CFTVqxIqSjezU5ijGOqg6/W/CaQs24b1DFOPiMq78TEfngWgzhPxPoIvyUezNXWu2njKbcDxstkx
ylg7pkAGn2wWBSH4cbV72ZW33hKJIKGJ6JtAbg0GGjORtXVVX/vvPlLt9NwlUG7pd8HBK9RrsRSV
sStkpOVjRWdM89EdGpnOOA0lVfaRHyvE2ExKVqDUzpmYlXgu8Z/X6GyLJL0O4yHSWak3gCWA/ThE
nt3m1iF3Pqy+vM2ejEVPnJzyzmwrjxIE9KMwWcGvh8U7i7TcxowQlmdtJAFEgZsSR/ntKFHIbjSE
0bazefYZhioaCakd8UvitAuycxiMb2Xlwgmvmc9gfpIIOSx56GAjEbdqsMEvYTBpZ8P3fH40huSG
/vkZ95uNoquzgn+k6pe7u0VrdJLCda59Q3QMfrxdNZiKdcPBvvgyL7A3XqcsxvEDJZRPDBVcYIvI
Z91MW/UkBvkiKkgXUEc2onzBn3TeJAe2OTg9F4XxixlTKpLSAnMApwJqUMyUI9G1tzLvt+8vEYdc
avRUn4/B7skZzg9CMrdn2MnVG05/VmRoO7feqi8lg1V1tVQCeiJG0ZhpRsLyEC2u8em0z09px7ag
nbpGPHJn8NhAhbaZ6qjUL4Utq2iQjhzlFT5PFZbEw4eW63NHWFHNGMKvdZIXL2QIUiXbTl04x7Kp
7XahRE+hb4KC7HLm/A6ha3kEIKdIgEWyioFjPJJmIzLVR21oNsodyDC4z2tNKtGYWQ6FUsOLPOKH
TvEfTJwZJ3V+gPueoFxlBGbyJEF/zdnTiSpw1yaTZNh3R0v8TysGj6XpFh3XCrScFPRHsbsKP1Cr
nRN2m4/aiZvuCvIT/F0XTrkAHqVAZYZYJh3haiCE0WjtPlN/mGKvT/ovAxpDe7NnlRpatSdjxPiO
FoJj5Nx8WDJEXZVB+SxH817LJTzGbzZNouscU+CmNQRpYYBflixpcfu4mTYC63H7ToX1dtOpS4IZ
aFD1SN90vgSUjzgpBHNUkrB5NGdLazrzUtPtyLiwBDmoJ/B+qQ+GNDsk+74faxbI58k9OLHJ4Lg5
obw3KuxHgZ0+BwGud4L4Hh2GKvnJwKc1ZBRoN32EiNQ5LC05nYKp4OCCu/X/Ex5F3Rpf04mA6QZh
cfIiXszGuEZbFcDUA+8kiuEM+eSwGW3Miszcn6Rceq2VmsrkDB386k7utDgjddEJ3mKspAIM2vfx
wrC6COAnRQz8EJJaSnndk+1FMtKkvLx7tfXdJRDGwEQSjKHQd5LDSpA8KmwYk6VkLy/olSk1qzZi
UrsGXw6z8UaL15YZq3ICkiEA7F194kLrkuRnoabunFsIXMPPMcbbcVeJbJiVwX5KH4aw3kKSEw0G
plZk0FSOTN6UF+T88XKxZF+qHG+IDqkhdijR8QAmLSNA49HFycYgvXTI5w2QVeptdtbnBb01/e8c
ulocNIbLx86KAUw/9K6C8iY/bGsBIwEBmcEXRb+3dwxpL8XFvLrs4GGIdTcZJRpXd8ZNtjcdGwLl
EKnU15B9AwoF+RjdcUXhfLqXlE7di8AJA1sUppFL+X9txSvrtvlIPmmqfOdvznxES04KKY6viFPM
43UdSGEipX1iZHn1Y4UT9gmPlYTMIIfNKjhjL6yGG3F62M1qpLHRL9eyfcS5YlF4VJLmZzlH/nfq
aex24/kbu27SDvA6JzuFquI09SHpIWFMEsh14OF4jTA5aftSbzdaBZf5q8wqCixL5tlDwfLbd8fn
DLKhtYXoGD9L79o4csfOfk4EHHWJLS94R427EHFOYZQ5YfSJgWJlwwQrFCocWhv/JLlDEWSxQA26
H7+kjWTH5xNc6C40Tpud/CaCWlQ/OK6N+BVY4niGznEIx3tJH6LwrLhfNbnUqmKWtgQ0tuEzzG/F
NNqexCa4GjLEAjbDVqSytLNyARchan6iIg920wxxNAHGBny2LzXMqQjCDZz2fmA629LYhvnonzvV
hktE1JPHASsJ8/xZi0Vakigp1LMYeiQkxzupsKMLsSemk3u7Y+odcUlmhh+jHnrUaua5U/CLFq2R
0CLrEO4V7eJYvPXJPSpg6BOyHg0VXVowbYNGhxg2N+4GoXZcUK6tyzrEImrSfAb79mLBDzmdDT4n
021gAeaiboaR6TKUxyYSXhpFkK7fMPdN47WUCmLcyapQ/4+LxPQDPsb9xympCYJPg9uVgBdaTxJG
bGLuFfAFBYUtGXiYoIGy3eiJs+6S+u5+ezKEcanzU1XK05WCnqvfg4wrDlh7QEyaSTBjWyZs5tl6
ZmE+2yN0Z5UqKbEFBzW2d0c9OWkw/d/Eu5IokrLtvzfJxQTbM2MDUvSqfySTeaKhJ8wA7huZ9C1m
V7qy1NW1hGo854VGuVx/AXqpWV4rDKai4Ft0CMXSK84r5CG2b6e5uGC4b0N/ZjrO/2PabnOI4LeW
ohru32X8Pm5toZK4DOKLRFSEpL0hsOGncoozw14ZtLZ2j2VwH5vfLMQr6LZH+aYnOjE3orrfCkkM
8FGB+USzaRgcsaQXOnxI1TrETjfvLIn5alwimmQBiAwAW/+iBUxp+W/pzxuqB6qKctSnbLJbyXiH
tHfDRaXXZ/lsI+oiXdCmTfzIG6e3dAJVvEBXFrzhsO8JkiNGb70D+jrGqwbHicR8VQi/wk0DjkbO
eWfjCCOdnZ4PGk9bEgauQqZEdjDzt3rdC3sj9rOIaycWGYRlmTaxSgO4fWNwcFYZpyvgXbvkuxf2
Q4V4GHXPSzFYfzILl28n3BjDTMNmsEJEKMfIWM2OEdpJQ24cjGmejM3DgRgbqqpoW+UBOGdxL70I
fBUAUxcljVCJoNdUi5oDsXmhctZJJcesunFemy9LQWoOKyt7BTs+lnYIpCr99HF+LQzZtDMZb9Hf
ApZ4ogdoGkvcdump3wsLsBH8jqbvXkZ+HXsgomUnljv7gfe0QDBbSbIMwNiH7sL00svUddej1BKN
jDAlX5iXl52lbVZQ0pttEn/QZ1/5i37qNe57bnR8itvZhf3sZPNW0ImM44ZRPfK5xlCaYLK3QCZJ
jmtz2eR8CSRuYDjgpulPMfBzxEp9gDig0TcX4gFljEavYy7Phrg4lJfe1APY/juLUjWJKtkda8oI
CAr6LTAQK0UM+CnmRMocHYqOI4/QrYFGFTZyodH0o+rdcnlbfTjfv3N5aO/oFK75hN/+ejCLjf/V
RKlG7EbyCn1e3daYfHmJnu4r1P9KB/Mq7M0WfXbAA7utLSDHMHOC2FiJPWPd649TBcWLOn9Ih65H
wMVsiUyqs3/XvtBEVrj8jKGyiUmhAPP5Z4tQ47pGDi/0K9EJ3ZHX9XIadmxpDueDkVuekjUK13ue
BSR4uysjWcq+PmIAg/Qsk1GeLEYMaakt7GAUNz5Tm2sBI1e5EGfE8H/OsJzixYG5IE6Umz11A2ub
mJ74tVQQU1fDfnBTTFXsDiqlT0ebHuIqiBquZ1HAkBjqQ8ah2LCSgCLd3N4RT1NnJqtdKj6ZmRvZ
NrRmx0yERkJbRadgZ5s2caJQRwr+pynrKYjPT85PGFrLHQpZLC2OAu09eczet2rj9H8gEnN4mzKW
Xnc5KuTW1DsxanXIp3ReeMFuzlpm+1+DgMGN4l8FG9SVEZqBcc5KTqM+YLRp0/QmrXNwGU+7S50T
UOw1LXV9c9KSbxb26yusgSUz4aUG/ozfEfTavgYQ2NVZEVS5dpGBU3qlZQiz3RJoXO3KrGooh/hw
M7jVO01Ob69sO32jvXzznOMQ0In3F62kBbaqrT64+EAbwGEqZNuaRqDc4TsxA0Ix0gMg9CCHrXth
1F3v9ZpuO8AsqnJp02/A3s1SUhAvd2EUv6h0Kh//znLqk78oSAYZ2uM07Q38UigyK5lIlR83EP8f
raE3aA2fxvtf5yl1duHjnhzjQi65Yo2lRkKOe+GcP9T/tbXJrIAmWH11DHI4RjtvufT7kPqbZzn3
0nBK+znnTaA5jJST0sP/odIcWSRL40RyYfdTB3YgHJOWhbVG01egRSt7eKSSgNZGHHnDSZPUKTnC
3Ii1J+pc61bgDkx4yuq4d2RxeorxpEGrrYL2hmGTQbPgJUFf8/gY7HYvPHo6nvzAlKrkdm2N+7oz
7b260j71Bje6fgLk9Xgk1W94sLVbQZ5CC6IEO1IgQ08t01nG8u92Kb+zG5YIVPREhrjAZqC9rcHr
FTrS4kY41owOZ9BWBHxQDFiNYuPGz4tkQODTAcOnWSDOEkDDoeUE2xymq06k2scl8dUKPUurr9qy
fCQrc8uFsxQdfEVr5hynhIDWG8xKDpUV/tPYhbMaNb3U8CWJjO3yCV6AcTJcHv2xK9HmGc08/Yym
qCiDLmOe0ROb6JJgASY1BjvAszEmaZKgeq78fGF39qXMtK3Gqqd2QjNRAel+s/SE4hx2jpsAd4io
KG7lmREK72KTq0ONA2fKgHHxhave3i/Q8Jrube3J9PSXbHfgZ6OU806rd4XMQf0GdaFIY2zmsyYj
dzkFyQLibooKixNRvfL00lRF4GyCxa+7kw54D7K2W+4pCQOOQGp1RpvlaZX5P1PQvh2QDC+6xdw/
F+X7pvvAaYr26NS8n3a5i3zAvBVLGRjX4100venvTI1z5CBFNkZVK9riVIaAQVVFm8wdOzxNjmI1
CYgU3GPWxUsLhfZYQU5xUTEVqOz7hp3f8sXZd6B06RATOtql8bPo2Ki+1V9Qj58GfgiRZMawACYo
aCuVqkTF/vGfyxeZdwlg11LhXf8IPLc4F/tSwReJEI0w0AqLUp2TBhF3wPpySs9Q70QZNx3wOlTa
6hjFuA5cSNp17RhdjU2SSRtWQ4Bj2wrMXLfs0ETUgue6tFjw1heqaGgTR+Qk9FD4yKVf9VtniDuL
cRYwq5BVAbaPxvW5SEzAs6m946uQaQV16y/IX58lxsiHonffqdxD2fqSvlFeh3Irwh5FMMtn+hXR
g5YrVdpC6c33fj7vf2+kZ9vTxAvo0nPSmzgQn+l3yHt3SXsdPqG6joWi9hutHAZMtVG5rfx+55TE
dZ50D5+4CJjgctxbaulUO4Yq7qlIK5wLy8RY5riBKOQIhUJ2eeMdwhyfR1SYaTS5fyfkmPKq9RVe
q1dyLV6lnft/Jis5FTufty8DNdvLnl3LIDHJOEHYDkfEMyYkMTd7/Q+jtzJW45XHtQJ2WUlFpqMd
2wTyl3FbKz+jRzFTNUcg89ml3jQv7weEHs7pnMcIo4lhkg/D8Xsu8ucKDit6YDMCffKwvY6AVzDb
brUqGeBcJQ+9boRA6fypj0+v4doIvHssZnswcmt3in82fR/VURc58a3H+6APGadyj07sngr5HquP
iv0agsy5la0BFuR2QYXnIINqeyhIzRCwhDIt+70kiRek25uTKLguV0y5Kwp7he2iKZAnQJB1trEP
wm/2y5rIkqDVuzt4vT5lDMGdtqbf6Fddn644vpY+DDBBhXLLVjmrF5hjP5IYQRzbHyuDEL+2NF1Y
H3luk5nlmXzTu8vYqtBviZY8iAHrdKi2j+mEnv/KyEEjMOXvXykTYHwYaK8PG1hRngcmOFI/GX+d
p9RJtIQ1kxgtulCdHg6OFwlOhRsg4rHME4ef1She1MPGeky7JpLU1npwV0wpFjAgd4mZuJ70kzax
v8+62bIGeDq5PsnfKWrKJCONtB0cgxAlTdq839LcGusdysRto9XMzZhO8CMP8fprBCRpUk2zirVW
5RXZwK8hF9SncqqM5Tdny6OGnjepNp73L101vm8pH6PsT5oE3ccBRvGnRdDFoiO9rn6NVHxhMSGC
D6xL84CyVvOdgATU/41Ru1iNhj5+uG4iC0SWItohDUwnk1kqbHzkqtS1HRtPvrnPYqdmNIlV+qJq
yy0whqgNPHQIOVOURvndpG7fMy6GKjxH9molMYARNqc4c8hXx7UUqP9hcsrEC03ePxKXeaQHpJ+2
dNfqvVM0yvMSf/Vk9Fgo1Z0oU/g8nt0Y9Mww1XpnZmOJxhFZU1blm5uq36DKlxB4RorfvDoX7plo
FMsIs1GZ3lnwJ+cpeTOquxY0fOulk06yFPAPEZyN4y3/V03Zfyqe183tCQPmp+Ui+c4lqxBjuulA
a9+TbSU2OTgakqGV0er8d48Z/yINIxKaG4wF77gYAwA6F2WZraW2Fl8HbeEXzqi2RiRQ7S6FW2qE
kplldQrbcUfeAiv1rcdQ7vi8D+ELvJzFkZ6V7ndgg35SYJ/O39tecubc2FSJwTpRV2stObtjfkF+
XA9kwY5AFFr/t6MbTKjO0TQRr3iAkZkJeKrE6FFjwNP4scW3WPMOey74xP3+3Org2urqMDO0mPJn
JkTXQIVZcHO2NXcxDmgLU2j/bSljEOw9Bcw+6uUG7ry/CXmqPP6tCFI0TxV64AcPn0nm5hn19PIQ
KbB24RX1ngPCwrYoY4wkpuFrbMGqbqmo6DhSZvY1oJMNpgiXI8sQLSE/lF4kwPHzHkAJgSQKyZnZ
eMYHgNhaFKSzYzmjHzYAlVPd4VnFgwRkQMJWjeamOwPFOVO3hMw09O9td8QCSXMROt8G0z0GvSNj
/y6irSePELWsDY9KIZ2EvORvcVLHmC0d0RDeMECZheT+CXjoLnec+uiy5bEgytKF+qbXLvGcDwCP
dUYuuI4Kha8i69rCGCd5+7Ei4Rc8TVYTm1U/gj2GuOb1N5RAlSM2W2NR6l8tyvJOImgE+7+8/I9w
JrMoPuPNhP2req7IzWCJa/2I4vF+wsgrWWvVPRa6JV5vDIWwvvc9g3iQv5dcQUF2aCdn5t9w7wXh
3xWNZ1osB7guLSLkRetHCYF92JTJPy2RcTDFimR4c1LjZT1rt75BCnQ0wWIaRyi77PZUUEaR0o15
khdnzJGeqo0S346Cp0i/blV/BfDRTxJLqvO9KgAr8r/difDEoJRbT1uCsLqYuyxDTJc5mlCms7cq
SX7zYdVhWLyE4oFgNd+509tg8Qa5Fxge8HB2LbhZanLnbo3p/w1DBomoCJXBBa/YEPmK61kr7YQS
7C0YfD4w8c5m3Ve22x5TyXow9teXZnGAIHHnpyyHWpMhRS9oUER/bPVCW5KSNIpWb0TiOGDdho0f
nFlPN3XigVk/EXdn4LA28j4uvRJMocbYZ0U2QX4XZwXoKW1FpicEE8xg/JYx0AYI4chffCQtTpSg
6KxxZ2IwbL1Iem7Usz0bJSijzl+AcDlK2SNDHvq7afUyeRYxKNsCBrlqMWjwMc0+DEhYCIPOd5P2
L+oo/sJMIfOt/NrKsi3uj5GaLCCtaCu+j+wnb0dSzrfw1cXdlKzZbTDFau1qBjwL2lb1jwBaOlet
IMsmCmZQ62z4X1zS6xM4nDPvBAwdnijkLE2VZXCG7FDEUbabBMRJ4XGsfB4bHixC7KYnxXOTPMIU
3GZYzsulYuHI5+hsKn2ULBdZgYFUdeY8aovLpLgZ6S6Se7pxkpyDtze/usKzJ1SgJlzI1Z9V2e3R
33WlVpEBtCQkCdELjkULigWfIzC1Tc0qOF3Qs6kK4iczK8ZS8gUdS8ru9LkHK+L4NuOGKIhNcGdT
OYvU+nA3wDCguNT7+UpqdNsuVXe8MLWa6faqZKynA0pO1Brbtk5sNR0hwOkvXjN52lPb4LSZ8tnJ
c1de8l8rMrB8q+q1mrQ9tqxmHBJ+y/LJ7ef56N+R+fEEMeHrMBo8vukovMKVK5t3Ox8kr/CvN5L4
EGDJR40JUphjBfCahwFNNMDQmccKyJr4M4c0UCQA7yKyqyCM2bvKYJAtxTy2huK89Y6beBBoZHad
f6kHf9TGZTUaafQGWFaAgxbI9EF2cJprZBDHuQ/59Sb0vJNU0fBzvB1ziBTDPRlAjw+Eao4Qycpl
e5pDs0I8VQEm2Q6dyYnR5QLhEESpd5yKozYCFPPF/Lur7FAaIu8L9VnkuR+0HrXz/6KMXu4RK+rv
2wOGPDFEc6dOqOtewTMRiN+XwC2pMHWMD2QVJbLP7g/bmzfAzn8UeQ6V9h2uLilzFhgX3C6u00X7
gh2dVjsG9OzIiEnNaMi2lcW2zAEAeS+NYJleukNqg16kV2Pe+SKnhCiyI2BqG0CqDTo7IvnyNiqA
vpst4OIK4qNv+sk4+zWQXU15wZyKeFne+TnPXLUvNn/a0+61vGe1YMz1v6BNFv32utOLjQs6QlWT
xVllNYudLpP7Im1LQ3Q01OFzI6YLkegtWALcr9eO2VrjL+Rl/7udHW6e+aWxVmt6Iveko6UVsiXq
Dl28GJ5c5V0THSNeE01WUq2P8eEhaxIXyr65mgoPsLt21wRWFJ0xT0281WmwaLiJmIjO/oxRWZqQ
D9kocULOjlwyy5K4piIkUCKsL3cg67isIpbtSfbhd7GQnFZpgieY83cRm+sT/Re0KRyx9JhUn4TB
/1zDjNXSmmISnuQW/JN/vMuccwzIasZMtm17OSR6sYydSnsdnJPCbrub0VBHHSiEvc2/QHHZdSsM
fPkZDuDtbF76AMfxwEOFVwg+6L09zX/zAon3gBnKVB31oof9yqD98HwMuyWQ1BneIPLXx86CmByr
AgbmXqpiIl8/kWBwE5B9jtA8Bhkd6m5SdDtUUmBMkYUjD5B6y0kTxBmJwku92RaMkjTdFfd5AET4
cyOHYhXHUdjhzi3naoJudoTGT/9rYLYbyEcczB7QiaI0EbUevVaFxz7ZanlaXnjcJ0C2pYP9WWaC
rsKQ2CCkzniNnCpdIbhZWcdYnEsm0e8XJZEX2I2icU2f47hP0wZvy3sLXHpgKVOKiWRQ4KFr5FAz
EypVmES31kbifM16gHgpUoUOcXG1GnNe8xVUO3AjCZOerWJhHMjZ3HDQ6wZk1mNNLVdpYPrqYOZx
UuIz6l4gIW2egZZ6mhAMsrZd5EThPAuSzmNz/i1KHmTulAUv97nq4PeI8LZihkArU5h9XDXvSycq
+VjF4CpnIaoTInsd2ySP0BJh1Ee4Jtvv4Hh6rNLljteeFkMk6wgTHelD6k9gMsYEPfRQHKzjoKMA
CtopuhyocXlDECawRRU9YP5YyWGahGuHpJP3L5FZRQN8I2himZgYf8WGT/IW1bpJdkTv0HjJK7I0
NtzYAzns32RRMsxjpFTJtQEtAahSmkomBECU9uUVCR4BroWuGsfHNveKT/mEXMAb8ypkSZ1sqJ8/
Bv69+nBNsnTTJ9BYpKfF5Bco4AD4+sbFZe0VTSPyCgQZ3wVngW2pV8jmJd8FmBIPOhVWIyWVJopi
gxiXxU47aRa9eHFqdYu3UHVNYGnqeEpasAkMVAk0GeB1JFioDeeZS54YAkmKr7Ps2eMSEbNqHmti
TiLCNQvslbJGOXGiQBDllOt9h1nzkNr1BmHi4r1EAhvx7E9gVtW512i037o2C+jsbDWy9cdkjxYm
kka+XZt0EJnT5oo+Rhi+tP0PNg4g0XyiE6tqPiT89wtqN+cKwaEZWkFrMGYG5MsfTABcdLjScP6A
OMnW4fhl2DeVmbmL21oCUAerqni9lJXACeVbqmji6CSy9Cin/4MUeV/fgmRn33xs+6DHA+Vk5vbz
atz22TVgGP8OKyW5NMoqrtiyEcT+z7TNy6NQlJkhyWb844uad88a7vVe09JQWsjxm8cReDDx8y4J
xcSudHj6jxJJOtK7vv7h1+YJMliijlezn/mDHyWMg2MexG5NFXcpxc5C7sjurzyiuFAgAZJndfSg
0z/lnBez44YbJBzxKwxGT8XYQfkDMFzbXnFp0N5WUHfHnsPU6Yza8ex3PgHW4TD4JZCSB6o5Z74k
gNbzgYk14kSIPR2IybfXGMtG4wIvFm2M7YZyPXoMJQJM4tAdpQyTadqxr46XDc2Zhayh6UtMjggL
rTEtWv+R8grXWXeukFaQYnvbLtDPXMbZfFeEoVgt4OFiym7mdONa2bi/QcNDa04Q4llAe78TdE83
9QK/PNVJpwvoegydwSZgKv7JFhbIJ3JtcwT8DU8MpzhZSctmX17/wGpgji9HTo9WCQIRlSw0aeyD
VDCAL3FbBo8JMeaeXyrVjDvCGw3chWxu+DJyoej3PTfFhFrcqKnoUfM6JVVHAYHmlgFaBaukjDci
DGDiU9plPSmYXl3zuW786T1fG0Bsqtn15K9DKoSNBcnZ4rEsv860ToSK5vEQ5YxDR9Ywlf0p08ER
0mwF4xBsYeeVITA/U9inmXyElwkQj8Aq+CUzuqVTy4p/bfpHBLOu8eOyEAVYSiMW6xY4hQDKw0a4
WwNwLhkzqz9p91TaDGqkt9qcuRlhBAaWmxwVX6p863a5LLWvHotTK7hP+ENRo6/frgtzd0vaieMv
EHyBxd6p811WaRRL6ujgJ+hrsZPzx80OOvu2Rv8+02vhaJ34um/XvtJ+TlrK+P8RQ0weeXE0++l0
ksuO42JSfgSvzgcRebrVXKOD8oitgFJ4P/4omnU52Jn22ycqPWDxtUlzpzOxpDCfKCduyRrNc/ev
zRWtpgSm9cu0mZNPwDGvQCtvBI3mY9LW4yhSpkb7lmcIljDtQ7usMGds5FKIPBuzYrL9Qe9CWOUX
20aewriG+B/BswcFPv6wtT1u8MO9N7zAMv7vO77cl+7wOfGzwV9clDKCkFVsPAjROknRexma9MoP
MVnJfdI1pJv4vIBnF1lOHd5XB6QKaj73fBzJhR3G+k8WGNkwqSI9WnVk430HYGSudp28uEZ+4gtw
g3OPPGHsSjM457Ev+kN0nAOAkijnkEQx5qV2/u672sl8I8V5xfRjgd/75lArNJCAIZX0123RXAqk
Ev+bnbfHUNxxYsvlwwgfz/O13u2gE7m0R+R/4qcByU+yQHTQPXscpOl9l8kXQ5ht/QOVBTusr+pi
X6jnWLw/nrvLAH68V6ToyFt4xkgwj+DEK8/7f46RF2bLy3Yip26J/MkA+Vf8cGRsmpe0wnA7XTKd
629QExMomwo371dSmyn4klry9VgV59tGYrH9+uI7wO4yP+vaC97q1wZBTwd+gppAGAo3vXj/EdS7
v6j0wG1Epun7WZhszS2u5PK6ndkmjFI3qW1g0M2FRmFn0evRnSLGFRQSLFUmCz9RMwr0Bk5lz1RU
KgjpncikYszkceVRq/gkDLuC7ojOOEKyOmgxbXb8K1KTfZd3eyQOoE0Mb6mEbA2OCTNon/l/PS7J
wtOeFHGw3r0pKLMhbkQLp6hzKnO1+t8qdFrXBJ9fr1MsBa9dFUIxsFdVCvoaI4byR/AjLHlc5oFz
TiYNGLrNLSfDStcEWyeneHX5nWcfIklmCs8KQhXlGVFGJBJ9jMam2Mi90xnAd+qH0ArrOV/SjK6+
T9dry7Q4JcuozjcvLpLAKHc2DrWyFXCagitc6s+7FrtraKfwZt1379ejOF46Ywu/uzgAwiW4x2RZ
azKoOfx349yJAcbNHoAVGhDP8bT74sp2qTtpo9KSF10AC6/ecSAGFtLJ/I5ilqsAPyCMAfG1kB44
hK4wMRliAGy8eFK4HMZKUY5jEQlVY0laIRPYFHCiy48kb0o1VrtJiEUVn+0XrRhR96Yk2NVdpjoA
/40nsW603kjp8zHaW9R4Mo15KylTOLd0LBNNI5tEOvXcu8tMHEwr+99gahuAyEsxdK87JNT1SEYo
axpPKFiVWPCJGYNswJQaVtWrd52N6eO9NiY1hGsfCqOqlgdA5go6oJI7WXQaR1ZEiw5jrHlkXvk9
RNTZl8wuA4Fr/hhiywv4Gsm16wPyB+ao0xfNpvNJ9mCw0L9NbxwOEpLpMmpSMKjAg3E7STmVoYuJ
jF3i0A+xipWSiBG1x/+VkOcR/gu33wEDaeJCE93WIhZFOwbtsrQkkO+iqpnKEJL5M6GRops6ebMW
i9K/ZsZguClObl4B3gAhx6oWjJKWrmdaXiCDZy3kIoia3q5tjZWZZkEK6IZjdcrBjHw6tceeloG3
6xLpBDGpkBHREGbNqfZfUxzQCjBS4euIx+Wb6yTWWoh+cqyfX3KfkIHsVFoS+USr787R72ZPhvCp
pU9eij1XDqs5ucfBx+lN9zkxztrO9XUJZcqMj/kZOkwMdipGgsead5rJbMph+jqi+ckoHd7E/LDr
rnVA1zy8z0C14EEyz+vbnO0iDtrNNanIkInzmARqdQv2GnA9SPcax+4tsJu3zIedk+mSiNf+edM9
SOvW7CtRaFanNfppxm5KXSfbyQfzcJR+VaoYk+SUdCocjAMoQGLulRnZxwBvqwwWUQQU1F57TEZJ
yAUixXMYiaDrs1EwumV2SVOHqs8L5LnKIVwSm9uRfXRxHopbB1MaXEd58UW1U6a8gOAt9aThxqCx
Y6/j14AmKJ3C/v5/d5yEm8pTimlpYDxVDYZPlJ6jgQc3FBhOJhqp1/QhuajhL16zzm/zM21OcnTH
Rs9o/4AE7XltOZo/xANFuRPW1moOgnPbFgbSK8MATKZlDx48Lsl82lTkSgzlF/BlfR4XM4J3AJoZ
VBe/3PaCKNDQWnxxlALP0ULfjG8+oUfRU5WLgTg8N8rEo3delNfkqH/Nm2aDrN/HUF/t9NvngduG
fqscK+Smv7aFhJOiigzGc322ZVY3OgyReEBbtK3efuyzCPe2gyAMbKpJ30sVq/u6SA60QW7ji75E
mLF5i/dZORc9yT6kAkc4MxMCJivZaHZVdccbMUp3UT5btoAny7gA8NPkJgIdTyvJSTrIeOZ8DAHe
E4FWFZJ1+6sRE/Y0OKOm6lpYaclyFyv+vU6cCrPjDjj/NH/jLu58Wz6qWpoFZoboWT3UWAyMnq0w
k3XFdnteRVrRJKTARXqddKiWXXOLg1VBAixMfDSMSU52614kVz753i40PbdKXpwCwqfLgC5BnAV/
Wb9G3S6FWlywlDc82FGN9TPgkLQrW4OOKDgeTiVw/zKPD73rdJ0Y0gV40IeGVD0KPBpZoYtcejFK
/nHqH7Pe5kkpKj75ydUrPnjmhk7+F95Ayfyaw9I3nukz2X4Bazx6YMfgOfWDEUcjE6nZfUe3qgrv
QJL9Zxk4F5GwJLSyAqjbC1buicLY7rp7wCJDex0xVwej6J2eCdnNlRnH66ev0yMYpU+zLkdyWwnz
vtCMOsdi6rAHn/Cx9lAQ8+BWIqe/eKgNCY41K2g7nTONTzXaHCsahpFqYlqMdW85HhxreUQXEgkV
SXngpK8KFKH19y0pCMVj06ddeGUujrmV4rkIVT3TmnsF28us7K3+MXHrN7jOwgw6dvtrvr2j/U+C
ibRxRnBIl6OFHDl61uV36inDU9TwtAF0lxEvnEf9l+Z3JdUROM6CKP280yQdpoeP2+ZX5lNCB57o
Hcm3wwtc10vvc7VRdjmCTBXNN3RezA2B0huN0ODXD4O3HOpSlyQAq37EwC3RXWt1SUtDdtDiyZKi
eCvyPTUIcW9q2w1I0FlrxtK/3ZLkCgF5IOU9QW8Dn1z4t4IjW5h1bp5PdEiWR89wGKp7llzOorZ2
N9OATuEDFvTRNlSwtquJiwEsSsKCoAovAhM5J72A3HS1PQiRpxpG7tmyxL1KlwzY50dwae4P9YAb
sG7YmCT+/y3z9v/yDbr7R2dnuBCh8XcpOY96exV6Lzr5gTnfkjDKHcWri2rb6NvDTP5zzHYIkmwn
odzQO0dujoh0TaOclXO9w2MSeeZQb1MogQfDa2e2ptoTqk0TIKorpWVa9tyqjRJp1zikpGjPOP3u
1YgowqrZ6ziirHQMgmaZXjQJK1hFgwA+N7ZA9rzHYjE7B9e8yRxnIch4whDuymNo08zYkxEXfUU2
iqa19vVbTr6FECQApGX8NJhUQoeSFOoYa4lqgZXoYRjYlTJK4/KYF4SU6OCX///EsEP48n/FYHXu
z5J/WDRq3Uq8NtOlXe8ERu3sO6Dl2iZW1EobMQ+lCBRZERwGyzz/LtMOB7QLJlzGroqsBAu7f8bV
KMRtIyHenmuGl4BEPxmDskRhkSwrEvB89l47g719qfEtAUOm3FMZldf9o4unrAUGrGNM569Vqndb
h+kxUYwNhIdsGYnXsGUWboFgaKg36//8ex8v5wYSYqz4Xa5lSB09ny1ZsmZptHWV459/ryQdt+sz
vUmrUTS3T1gP4M2gend6265tL56mqQgf0OFwDh2kyHv09mwYuVyJWNJGinxcJVfP04hDbsQSrPFH
RghdCwsy+VTRybk6fK2GkUjGZFie6eHuaywrYay4ffDXyldzY8LiHGuqEfJn7RgzwXiYaQz76Mgb
YNtOycq3y24RVSsbnkslEc0toiMuXDMr2/EvYBsvSPoOrhehhAtmPcQkCdrLjjlpQmyRa8vrYjFT
yfabG0kqego7rTRYOYUithIn8CWRiL9OboS3Ey5vCJKbE3iszF9G6pl+U9rFq92svaS0AOi+1EPM
fLqg8JDn4nwaZRyGv/8OBR7QgOMD5QL5bPKb9y7L50T8lM8LsJAzP8Suu7p3JEJG7lXS4+OjYFVD
KQMIctpxEIT6l2HmoqSuzez+9ZuQkWGVqWSZhZGDFpdoqMIwV0WIB12FJD/NNGvn4/WYFXu5Qcq+
q4cyVfkM8AaiS4tJ/ITPgH7e1GqzjqTO+2ThmKITUmMUWc3nyhfRn848LwMipO5Rv+pVc08Wftay
HiFn/zPe3mXzZmC7UMeKPXJgkz1LE5DJ17V7CVi+odDCjdecqFmpnOQLu1K+ZBE5Iw8ITfIMaRhG
M/OxwL65naV9uUxaFo/RwnCR+YdLWhkNWIxWwFPZMqdGSCAqlTU41iuk0Ye7MxoOHqrHTrp0QLip
RPsSUaEJRz5sdZyC1qIaEtimhx8YsriRfQ9P1lk/+Dq/PtzzLoHZO+rtZwyhjjKPCKgoffVBcuME
I4pt0waNjJnbfgtJB5+YimeoDmHrPyFhI43anXFQ5azxdEMQ6o4pqGsUUs0mJtidGNnOSpkT1XNk
VcOwZ7uMzYdl4oTfsNYfecb+VefkF0i+PpkBddCAJGF3jwbTSXFN4UO42PJKt6pK3UXuFHB3AzYR
oot0+gdIasIgizDv24/okoVizQRc9A6w+9kA7SXdE3aMRd1oQrUKyIjc7UopuqRqBqjd2bn8Rjlz
jfBnfHtLXWjJfUV0WmokVlYyQ1uDQDlsrz3EqkhmXcXcdzEOZZaiCd02ZEX+48od23svFXC1HrCi
MB6FMpl2poHXr2XK5oz/JUnBfkh6V8N90/deLtrMvRLjI2jdZNCoR0KzH5PbmhxvBhhdd0c/pbiw
wBz5obIIbMFscac4rF5k9jx53RzmP4mIKvwxBqqDE+GoNZiI6k7AGiFj10nJ3P46LCDe446yVQyq
gyvcF7J1/qyXMPWZkmci1ksNAB2XLx3h1OornQYvWVulAd+ptNP7bZHghbwN//4fxmXE/q7/t91a
VEfcasb5khOBr++sGZrVQzJ7B7Srk9p44VbPebVCyyo1/1g3zFjo74f7gQY5XHYOK7Cj6hu4y4Qz
19stlVURX+hq68e5oST2m1oqrzadj/xgYl0KjRvuwH9IKqGh4EWd7TZdNyM5cmnN0lbd9KCYFqT6
n/gJxyt3oQXrmmJJrti8jQ0VQvl1DAgK+CKAIBfsj8goP3uVALrGTG1LNG+CKTp2+/4RKVEWfLLn
i7fM/KeD/gVM4A63IZzz37us8lBu4hYMi1DxMI7qz3hdQcrEP6MeJpt0dfaUe4RaZ8+pfQ5rCf8+
+0Tz/xdOQJaBLf78s/aUQTJnzm8wgszzM26PQqQ4vaDlTqnEeyK+XYwSYTjfmbZmrO4uC59fNGgc
wCp+LP+4gBlwmz3DPCUPSQBd98/17DTbsZHY0GYuyTSjr0Os3cK81SZiF7tnreqrGTNQljoaBZjt
hkeDx6G0e2YwfjL0p2BlO7CeCwGAhiHxlXr38Zphx/UuopJsM/jXsEjDsbw7+h4gp+mrD0oJ7NFS
Xx46rJXF8xMAs6o+blMo86018omR8HYY1494j4oDVcoTakMEJhmP/g/7SaXMgCX4l0+y5+I6gH7K
oCylQNTwMUbjFalFxTjs5mdHdmboTTvjZJOGjavn0qD/nysQ5qiKQ4lcAV1H8f00kfyP6nrzhzOs
iY8iMV+sQ8Sa/rdj1DJKDcpusRtp5Og+C3jAYeTfEAyZyaAElx6mdYWKQVN/WHnGiSeBh9sTITKA
AvUAweOOxyW1HMmOeUe8XSzJt9RAG02uW8gpJuHqJBjii2LkT/yk8T8GFjj5gGOJDsHj7o4uJfi4
t0GVZV+msJ+8L+ZlxoDXDHNnR/YwMJmsU/LFC1Ywj6UNqjHNulMs2pucRqr0QqCOm23vtw4mxf6l
fWW8YB+FBwgmEKrXHPAK3jOPNwacb/burMykb94Uod+o/tmDpGhoSH4MbbJj57rBU/ylecQdf6Xi
FIOfLBW8H/HUevIJpaXNUPsgoQphjedQRpIsEDhm0Hs33BUTdZgQbXklTK8ABiLBkD98M3CgNtZR
ntgpG10pCOFzZg5cruoXOZU+voF/VFSe20eBFAtckhBfOEVXa7Wgqy/Id63oESjKv4V0VU/nl6RC
4dYETtiRasnx67n6Q5pZCKYsoNDFnts5ZBrl+AxYHHnPT/Xiy7VdX09SlVcqXOtsr3obAhsXatUx
9Ioy/q01CTccwi5bNO5p+gD4dATdomGLc+RYtdG8AAQgQZfR1s/omkm1SglLKrfTy8tzslZyU+iJ
AvoUE6zXrEA3nxUR2JZjWLRboVegd0gIWbkjkl+wsZ2yKBayEurHkU0ZzokCK2ZGSwjKWlHAuuGw
izFbla+bive6wlOXkVGin+sFOit87NndsNJs3hyijvLEmys7q54Q44tgRAFFYUgXNf7SvsAqLjhl
Eteyy8slhst4fZEQHObIQnLpoaXD5nxBEz8H6XkJNyg7CpXz2WBKhd04ncdDSIC4CmlxbjCTn0pv
2AaFqjtuh1fq4fcPIrlDEM42f9umU5MsazTusLpbISVwXhSSHYRx6j/ItnkSE4HecXaeEe8T8Ldb
qAAEUWZW8NQdnDI26J1jx/wDTx5AKqD0dxUsAL/iP8tJaoSAVc4o87XxuOgjGjhGZRKcwXkgsNi4
yPYhvfclSy4wzf+qFwGl1UvCQ6UvpxaE+/jDwmwnq14aRDuZeYhxQg+6x3V18mz63HTKo0XUKokC
0Cqht0RmFsnQCD0+VdWxeSL89TpYBA6MthYHvnIb7LK2Afzla6HmkjSBGPaZIGnW59ak3H+jETzV
ioCKFmcxeVVgXmHN2cZe0lheQDNzfWKAJ1ZaJ87dduTSxLt7PnrzO5ehwyseeB+htXCm8ZdNRwAH
qiZpRDSwZsjmgcsDsy+DJgQcUnqNmqj+R4LTKjmxt4YHvYp3DnxdPLP5NKCAWhKWvwp0vhFYNIHw
0PMmNKVxpyMV82Gyz2sqvPDkwP7ObzYKDjicQHHrwErcgLlaOWqMwe03ulhIu/9AoyhCpBO3Yd1m
MFiAXhZ7V0nWtOZL51JJKb0q7zPLhi30YQEZyyMOIDrfbLS2f+KjTLD+v+EjTxCws++tX+TyNAv6
hsZ3KNw6WsOQuLW7EFek4iokjTBeeak7VQ+q9fH8thjChr9VTb/8W3ESMAN7g0tuP1FVIW7F2fK0
fiMIlqTL/1x80Q7OL8TBOpDMhv0mP5HmnpWpULp0wZ/jUxDouq7ZUE/cjyOKTUnRdG7UWo2Gl6OF
yzvE1ehfBAkAlQwfHgIDvcGX/GLdT1yJliJBl2ebzskR7z0PfZQBZgOX/EFnM/DpNs/W3Bsb8mtP
PTrzY6Dp49QmPAPtMkcV/8yJdRA8vedk7jScNlqSivJ0fjUMQJQ9sHMr/Jtn+jcC6FNMk5lnsmiS
fanFHe/+kjYdUAKxsxXeLJoT7EloaEDFYBHeB+nh5Oeqdsl8c/aZ0ILX6LpkC5YM2NQJ16FfjCHU
GHzPkz+lDfXK7gvluiTe2W58znTPWg2nIYJFvcpwfKxvFFhFApTt67n5FdxLxcqNbetFeefzJi+T
pDEPZ8q9dFWkOlux87bfO3r2OZHxxDBT4qrpYZBCxfT9Jrm2uaxXTb77SSlYnaID3tWAkV/sHzK8
MgV3EwrPlnJqYrNbsTpj1ccl9Eyk6xUX4PjWvhZXIQMYzZlvzpyAjTrfh2b0MPV5tjSmdPg2l3e6
eoS18Bx0ZpidAoRw+44uUdjMG63NK04EpmiPWukQkztBeaOFaLSDDuuZtXF3cH+nihlvip0fBCqN
1AxOlc55wuS8YCdOrDlHdlECwGPrjoUoeMP3kLZFMP7ZlEfBR0iTke0xq5DsanL84EWttrNZcxxD
E2K+pfArzBGAzxL02vzlmplwwWNwpBuagrwnqQkjN8hsg6KJ0XYoO9L8KB2+9/dqcNbXBs9sUAWN
YLXEtuK9yxvwome8YzXBYQEI4t1KHxR+bAILk11C9j4BGvZcUAvNuYCa7svSzH88Kqd1q9fEOpwT
t8guXxR1fPU/zanLqM6P2dsiLcepSurhaRNvTaA7DmZn4QiexeAC5xP/NSbYkXXX0jk+3vTjYyNj
eMdchcnyGU0W1cQlEJbNRW6I+BcTKS8QQotklwHbUE25DKkPgYSdLVD5gmBPd+T9Q/wFcl7j4WxM
WT/bPE/s3y5PLwwwqzitNnbWp+1YQDdSVeL2TZnTtjxutKUrhJnIGJYv+MiNj/P6RQYH//M3YzR2
LdbVvX4tU9dYQmUMQjVaJX4+WEa99Hur6afcajL+Gfno54Eha33LX9moWIb7/egrvZ3O3gSLEDOU
YwoiHzxoC/xvxGMoOUtfIJ4dSp3aZePPXSMbRw0bXrt/A+gaWTAswuf6OQ8qxCIWlgHJjSJBjLMF
JYATUz+MbfIVlA11iLyw11bskFOm07O/Om/nZVtLzu/b/If+SSVFmVU0OXe07/NQPQfaoL4TGq0p
o7wwPOC1oM1H2FB0bDg0L1eq22B/pinq6N5KSzOGJ61xv5VhzeqNHOlmUXZh3aJfjJz8Lf8uEBKn
CkLSZGVmJhVf8Vz7bRyJ3jB1Lqd+ZFVZfjFRKUQ37ZfQnNDWvQV6OLwlAYVhXQ6LT2MycNT3uqMu
rn1emS7dRGM+MjFAYLmN1xvQkmQN9viAZN3Bqq4n/mjNl/wco/vgPZeouTFVvIZa/MWzB4qEK2jg
fryjTWniDJeO6qvcVu3S0DJDhRd5+RJHnkB0rgbbjHhVpS9hMOaGyYjDDkDSuyeNa3u4pcolzgYK
CXc381n8SKnwZeVAy+WiFhLDKfVK7nLqLPtP0Wh5N4i/bVOR6peMHmjZTBcyIvgAvon53RX3kPb0
+FcgUm0t7OQXY+uAaOCB6Z9upse27E6p27dA2Xw2lJ+hZK9Jy2AD2x5hkElxftmGG7W7IpsIHm1N
kmEdwfcVUDqNEBsDvU2dS3/O7R9cFBBBGNnF93mLt086ZdvCQwIJJoteXClFmLaqeuYAPb5wi6bm
0kyCU9O08iGfWvQqfRkp7vzxvgpzO8+3NOFcJt1qYcq8qrGtBHWcw/YLxwUuOZl2dDM7+ihKLyEi
fE8C7JTgfqCBD65lkQsaAaMGwI/tMnh2e1l4/EiAoL9MmY5E727caWBn6+ncfYg3yJ11OfF/g0MH
U0+uwHKnD+C9rKT/wO15MnmEaAsobNvjn5z9+JTtIG1ndlxcEJhFWw+18k1Zoht1ZPV+hES4vIHi
rwT8+I9HEhEA6wF5YoNjKz8tjf+GRluvupNlDZ9Mkaem4JMcuMepvOF2o49TxqQ5TlJcexTm1N9q
PO7hzmW1Mhx7qRiw1oHyUewIQ2Z5A2NyyxfdyAUUqLlIzRP5fHfkmHjsOsDbo5CcLLXkmSnZa9l7
ANgR9rCdzUger7p9eCuZf0SLaGD74AsYFRDxTwiGUDvWG5Jd2wOQiwsD21566W1fLp9G1u0gJjJ1
gnP2L2GvxOiffzPDZydz8LRq/v8I+hPUHaGZf2LfXOBvsorDCdOQyHnPZxeGVRgX0UdqsQsRxcg2
PrBk56u1hhhUzPcOUWlN1/PdamVJeSCKScgAVP+qJ0AOozCP5PIhCvFhw9vR5rcBHLSDWz4EJkxW
MhyfHtLDjGPSMx6rW7eC1rtG02U2ulIToHOqkQIC9nXso0BGF6E3VRcCbrhfAOUtabbOV5UClx8k
Nk1WXGvLayG71rf8w7IJJ2rI+3oxPXui7gg/ydzXkz+OjaW3FjROWsOIZiEiihEGkYd1l15JVKzB
FAesfulfcjudBozQfBlVoTPfmQaCcttkrvHZjfjUZbTNmwyrK0JWWGULzJDxDLoXV56u8fvIotxl
FMF6rf3v5RL1ryRPCiHeoAP1TesthfGF0UbEQvva/o3AD6xDuGu71RhUZ5uO5mGR3kb/OW33Gp2r
YKKmUPt+9+cc6tdUuf3ExlQj5tgq7L41OiALrkk8A+iH5HVvRmZDRvefmynXpkSxQh4WMECLTr/J
B8oNnDDGtpkGtHdUHW/1LW8gqoIyt6G818Pvi8/8uCJOKb8ak/vRI7ECjGHItYiAXa8W55caO0pj
8T4yRQCoNE0bTXSdb0EorFBBpM9+MbkXNZKOhpHSzWTq4C6l+Y3yrS3VbOQhrPLCZpmFWa+pJumc
qIGYOst3quZJaHjGie3ct31W4lrQOh7Py7iVvpIKIftU/pzG+SvCovXRKV0QbCf8NMYOXse7I9YM
oed5YE1Jl6FMc5mKGnI9PbAc6IURggIFc9d98wgzSU5RAWMUjEB6FSPa4l4CgYI/lxHMP1CuzuCk
iA0yDeALAR0U7lTaiO3zCccKTLUJOVo4L742TLrmk3xDqIwwUzW3FRwErgBWCUc6LDo6BG3/ed+t
lLPJsQH8QV0nlvYdSc7f3B12LPBnmEp+eJuAFtO+xPdJ55F2FBeZIHt9sAJv526E1p2jahqT+V4F
1nQrlmTWTYiQalnfPd78mwTtdyWYA68uCB9awokc+uLtGY2O/KAYTORnzDbV7Q2+Sdq8nH3g6Jk3
X/dKpw6NOphXzNSUCe9l7wS2t7cJiSzrP58D67BIa5SXJJE98Fs8x+GDh+zmyb8D1neh6ND9ZdHA
JtsL2nphiPOny13ryRT2J8OZ42twurTAURqe6/peNsEjxPdFBJVgC/hkDTuNHOqW4Htg0+v1NnwN
lCw3n0rrRR1zGfSwt59LAMRj1YW/Ks+rDPIBahrYMZp+f3UDaQ9m1UYF0Pjq4/TCdhi+u8UyGoQH
rytmi9eCFEopXrG92o5lSlg5hqH2HkQYh21dGb6WvbPnMgUlfs5+vNShqOKhmSFL8rWfDzZnOoJ2
qt3nxoW7Y4IckXhVYpEdUy+m1P1fEzn1mjoBwzZLbuT+vYzamNJhNk9XxZdeGjVEgqsmPotP8yJz
/uC83YoM+eHCTVFsovnB80sLdMd5n28euDE4E3VrW7u9LkC+jwD+NAuDO+OmInewTcXgFgJ+EYnP
YUQ+IvuyYAumO4wtMmcjoNQzbjsQfCCzDBFhJZnnjfaPXBpmpEqDcVNwzwxhcgIFkwn478Xr5QMs
rb9ub9xVfwNZ/bnA2Mo4LvR06v99bIIQLp2YjLl42CxL08waftAa181HO45VZNUFs2mR/yxVd52L
OjSl2/Il1QDuhcey4DjRrOBO59UqfO7rJolSRZ+Zh7Y0OgOpNZa+y3ToiCiK/DfNMiHi18hDAHRd
OBWwvMWgD7wVvWryE0jxX2pkUdsNwrAWmz+UaEBawsVsyFGF9JfuP4xB7uH8yrOjNnD3TNbpHT5J
19FVuEWGfcTGYVZGiMLZDrdIEHiASTQO/cwpf8UqsEPuqmXnWTQIvxbxidbxLm/RxieR86j42pCc
18mr8aXj/Auqzz3H+6NhJ1hxLdvBjBF1s6MAABbrzF9mZtUsESaUT0Ll/5K7vzBJgYk8T1AlfTYc
Mwqu/XIMi1KUQaGJ7byDZExkOvVM1vc5AVHihahHbNnAk0JoJf4jG8i0YrkZNYxI5JNM3wlozRD/
RX1XYsreBqj4yP9qkF7NzgLXxf9RI44nqJE8Eksi6ZoGTW2xvgHCHojMkwLgH3k4Fcxt0p6M0trJ
qy6OWsdM9pmPsQqWq4KXAbPTXKpJyB0he40IuT4m61Po5hU5AT8WYQFTeSY9SNdclp5wTaKRNG0C
cQus3u5NsgxSoVjZla1UHUrB0WJs7wBuLrf42vRoe6HqBB2rv9Y2VF/ntI0TMlYTgFesKNEG2wnz
h6mgONBu8NKawm+gfeCVcMHLyuIWPwjpm4DgjUdrrrNVt0LuqbouhAagTwUJGqm8JjVbkcnWpMu8
ux2htJUKDsKFZ9ervmr8oTwIniLSNp9w36li3WWKlyx+Ui8RMAAoqNBs5na/7Y5wOHaR3nLNsD5m
qqfMTBmBpsG9v8ANv2TofvXyYja9RaqwE6d3DcGc04k4Go9J829wpR6dQA8USARuz0p2QsrAEiNR
rrvlPpFNHex+pwxnKqRyZ+Kq+62VYRCVSAXlFvb513FdVLr4bi6rpzNwUumaNtMgTRSVPG7/MOrL
6rt548M4zRy44L6RbfoFc4INQm333nDidNI1Nq2dhtka1xhgz4FWympc8vCWnXCvML80dPoLFFJa
IAI+gHlwKFTrmY0UUSQAP3Dv0O4UytFM00Yfd/h95BtiA0vMp3wKOVVXnjpx+OJg0ISfy+x85G7g
EpT604MvEUP2cSbRV03hYFa01GOgIKlchCU1BcYXNjQ1HT/gqh2CAAyQOIITauHjrm3Uwbobxs7e
w4UKoj0UuQdc1VaEArjWLEWpA+M2aQi9jng1YpTJ59PtJggES44tP4gSyT2NvxLEwksUc7480vgz
2OokfYelt0Gd/9vi9zi8XV/3+fa9JfbB5rGAioH4LyJ0vf0Fz+/vL41binG7HnmDrTtDotIE5jWE
ZdiBdShOdfBAZKoJyGA6ZQGKvT3bnEXUNzX+Q7Dn5ymshyrtY7NSH5aNX237TuGNbLb1hEhRhGK+
8cyQtv0W2Xv8YmrDyaA2XbcMy4WlUpA4DrcPYtjiYVZRCDjgxKCHlloJ4A0P+Y9xXYyHWpX/GLGW
P44axsWswtf2ujZxKl0ALYf7kN+ZxdrF8Om4R1aHF+oXlOWgnTl5KVNSkRPDMQV5C4Xy4xIX0dpn
IE3amK+/ylsRv0coqTnFnLDYGrxvt9nhZ/Bpdpf25IZVEg0DdvsU/DvD7hBqrNS43FW3/WFqXjgw
V49C7xV3quWOMehnGB0qlljf7qNXisEYTzRFZN+DhNmtg4XEdiDQYfy07IAJF1pbjqycvo7Ssw/p
uI6cc1Jtx+Y2BINzNRSW2lh6jEO46O6xDV0uKT50SUUDuKsIN8tRR41JVsijdfG44o8jpEJzC6xd
7qKyUUNAcpmrBoagWqSHPZHPHcScxa4dHy6ARlsVAmo8PB2pT/5Cb9Rih12b/F7NwqABYDELuqjW
ZnMrava5bexVVb9BVGWQy0oTy4TRojsL1vLd9TENL6Lb9n/fn9L+Mzd88t5mAku3mK4hnRePHcxA
DSio7IMA8Tu01wTbhGoy20TQbrW2X+RjLVytxVqqDiJYvWkd2N2E5noDDbuBQU1+YwdBdNTAJoBm
dl+C0h8TPGXPmhoWe/BysVwlpMxSUsyF1eTFprDjqsjTgKnndGkGVfFRm3TkCdUn8Ogwr3t50hAs
cAej3+tb1DHcPHOTjmlCbMqRIREIt+GfrsxE8YzaKexNpT37cmnP9edOyemfFUSXnySEMRKegvbj
yWsRYx3xqQ8HDq1qf4YZNlGYQUvbZ7bBuQhWEKWU52ayucx9MOuhvXJ/6BMadtzeIWlMf2n4Rbru
tJPKlO1wKVeq6lZPyzMW8d2ZhmuwwsDgvGBnk6Oi5ZsmaqHRoiawqAVKbxi5muWH603ocWO7PYKM
rIyfdk2/vdxiqqetHnIwaxlvWOeVmSGPOeUr+XGXtKQPuBZpWSD5os2ZEtAzilUDQbsdNbv8SVqc
yO/Ffce6YO4/ucNK/wqO/sCwW/HHEI2Ay+67aP6DoUF0gp9oS4L+9Ora8H/Mp/MMGNU3KuHPpsBY
SxhhQ70zngpzFg/Ph5UuVVA0lbavl7BaIhtsgKf233XJUj4M5PvCsM/1+nIDv32NYbQEYKfYO51r
K328cbOPFw2fHqJbGZmFXvY5wGP5C7yzHtAH+b3wP2iaxhh2r5L6885uh8jupDibxbxNZVENL3tI
YqBp5C0E8zAQ2dy8S6i1FWV5asi/vHEsKiHVn4y4vurAMX4Pd4Me84TFenb6KfyE1Yhy4BaFJgz7
rF+/V//NNZ866dU0EAxb0sRoug59oXKCbOndxfDMutabrOx1eWGS9xSU6Kl3R2rn+9jvg4FD9ukr
S8PkksUUtZSxTgz9gz95noZ4cpR9kqBnqj+GGHVQBrMrPNpBQ1wkmUtTsJEjiPZ/4tercv98eglj
0mh65RT9z2TAC7J3Y69J8DytKHD/yecg601PKLg4P5UJwjmjhInYglddmw+1phV46WLUvt+5m18G
L7+MchYUuWbOYx2xlzzCguTq4kAQ7nlSBSGeojmvAayTpjf6jUrFWPK85tdrL+4uF1X/50+OAi5m
aD/xI/ScROLDKmwO6xqQx8XRsX2ODZS5QWkEegZDDi3P9nGB8AbE4c4aR9q7ss2cvXbntVe9r6Fe
lH9BOmDOyboJiExNEmYL4RQDWXplW3uU+dEjagEFphgmKDrO0Te+il7XRt7zvMRXFw9TiiSdIGEG
12IqK7Wkem2OL2ucQ4YlaFor/oXgthWHl2hXBuae/SPCFyiUZDLGSyFeaaYdNjLOUPqaUUG4LOhE
cqNQVo3hooFyNvcQkKZCozo+AxuAC6JyxZrpMEpmrc4OW3PLCTfKcb3EqrZG2EFiK1RtkNuHlJQe
VhxJT4s0jU5tymLqc3Ij+MLaiEQtEl2v2W03nox6i/I5D6GY1qLyiO1ZFhsdwjDoEw56e5cWwB7i
sqB2bZpvWGIzFwV9t80TdrPmN3xNi+0k8+1+kncRgh5zFzAYeLVdzkqzRNZCyYyTHHPN3cGMoFL3
i2aRohBeiEvR593sg19o4+GKhvbeXv6974DUd7f8FFsE8KSFe9KcuJ9FIzTWviqQQSMKw3/AUiKD
OvXfSWnkuRJh+Jcgs7VM5eiOivxP5PAe4pzPtn52olDYog0NztKcd97c0vOPnFmZ4rMnzZ78Nw2c
XLoA/lRUu2jHRsYkACi7LiaALgm2Yp8Me62queOt6wrKdoues5JYHhnzl9/060V+/jDBUTsOTALF
6fFSIAEU2NRqdEE0GZytuh92beJQzSbqZKD1Fc4rGQ4MbVN880KZ+FLH3wpLjDehIHgBs4ceVTAa
fZIDU8k28IALzzGCRG+E7nLDgFTjQoOXt8BEi1r/BcDz+U3JZLc8Jujdvp0B5IRXkJtx3eZ1a49Z
E26WjU/1DNn6QVjTxT0x5HobqAHraKFDYtAASI6t3B73Q7qmhBlTVbI2YLM0sW5JdxPi7yM0ABRp
899Vv2ZUoJ7b3CeJnlubvzRbwiOTvuc8lYucKK8MHyHz/UKisUtJPvdFs3Gpjdw34AYmshxQicG8
82nLl9SdBZA1kndPI+f73gwXUBvP+FFXA0Eyzgy0Slv0ADFrfUJYxMoBWwmudxLtIYFZxji6YOgs
CfDH+H1ihf0MlyNTip2/kiSKjmhHM7ZwXg06bvfs8OyROxZGU5lr9dilgKJRK+zZauwQgoqcNroV
gD3UxhTngEaVdlKP7AkMN5qvMgDmequFDwCFXn4hVHD5bpbXYKQ5nM8QJOgWPqZt1E7pDmf903Qx
798cn9Hj+8vLd/GGTs+sldbLFjIWMKsRe6Enrb2zLpr4pzkYT6AoEJqQmzVOFw/x0YlqWQdVXasm
mEjnPW3A/ioZklamAED5Q4hJMQ6ze7DJnYcr+lw6sbLUBrO6Hwv0KWIkRz/fGNLil2BFBlti46Oq
KpI98vku2WHPm3ll9Wzx2VhGn7h1IyemxHQFVGKX5mlA70O4O+ros+zTbF6/BeQbJYACkT4gP3J0
i1QPF5TJbv2VJPRjmv/9oBhlZFySeSYqnQL70g+X2M3ibkqYXGD2DATTYr46vX8EK4ifF1ZPRPaa
CfEAtGxt2ft0/e+NowwTmpLMI9DF70uqSCNqqLLlE11CQgOh7QrgiknnEIr+z38auCpGSePLPuM1
WpSDxMQfSUiUTurV3s6CHpwVA+24Yw8Ac0lrsJhh5Pzioy/+UO/tilVlx32AEbGj0QLjoNZeAjxZ
QKikBOxhMmHjOzvuca2pOVAhMUBgiye8udEYB5Zaz7ZbHW+7mgwlcaxud5fvUMw8HxpeeR3VGdjA
BA2/GbwfGGwth5eN8S/qGKj1fMAHaCYFrg3fMBdRxzudwJC8kZ+NRBwaq04+VaXxIwQ0+EMNPUlh
BV7ySk9UG6qu5kGIBPuwOoNJa5nUcYptPPMEYpJn5LlTR0onEoqEmCrKz+AgfB9t+sWlJJICZBpQ
eTqa4jf5CwIzdXvgMBc8TblVYuKVBIVmNpdgtnQPyT5LzLHWTvlPJVMZKFEV5yRW5PxHMU5S7pAd
PxjX3+n8xM+akaw0OT5U5eUMzz0zxx4nKLg1K1ys1YcbG7uDVCSI8RbXxpqf6g7acgk5Y+zk3hGZ
Ga3bUiQMcKLshWEqZyEzdHvAXIe/6+4blREkKYkYZ5FjLch7gD0j3uIBrDDmQfhLv+jX0+EDA5uu
UvJtf7f0JDlB0cF7nzbfVHPEL5s89324BRD5GWbKogIQFxxc2wYw0m5jfWh1JHdqcMOW4wcEu9Dl
8slLxDxxJl9LY5QOMJTUBYKK/lre/g89s7FzAlzihqShlflEoAlw0hC9lR4fWmbi6dLYgxdN6YV2
nTGqOlnretvb2Gmvc1CryIw7XxGIdoQ+IX8ERRPwRpgkAdVEZgkO2tBagcPAN3KOyfcc6sT2aLpr
ZE6fMxrOWsSLTeZFZ0DFWJstnElux0je+g7GHdOpOgID0SyIPL0xCAiNhLlmqLUDx08gn24/Laxh
8iq6uHjOHjxZNEKpFUksTH7w1YuC5lX/YN/FAchphY2/eGhGb4EB7YZHmPnmLXI7QTKVIvNLto11
oainD92Z4z+0lh/OiMZTvx+xrO4YcUCLLn4jEYAJ10YNEbBGsJdrs7gFuGtVbKIrXCLVYgMxCWlR
m6kds3MfV77+61vRMqNIr5vn7f/acpVY8tOLwM+208qyX4o60T0ojvCbjvZWcDTOnyAf1qKAR0K/
ZRNFXECiVgh6fVAmDjr2pmF7GB4aWZogWnL3e6kE8Cd25glqC0nVKzzEWEcYC62MF5V4kcGYLg3i
o+nK/lXGByMrGf7Nw7/jiypA8QnHvi5HTN3kPRsMVtL7p02qX7o7X6DnJsONdWA4SS0vsk9IDyME
02OeFcr8NHw+xQXwrwhSLhWjkjX1f4UP5IGbmsmwDwUdSQNTSqHXCm/yXSWWnF/+EN44+L/njKzS
YD8o8JkKOC1irVgHO9b6Y9XZE/T4alYE4oshBuEdPbGgVb60vt6xdPeRc0WWCAT2glIWwGxv0MTj
feAxCuWZiGHDB3ZjbmFMmcwaLRJXBN7RMwdivXCOq7ACRX192wpeMQ2Up19E8btxGLCQ0colvimS
LPBOgZ4BHnvaGO0ZvOf5kCTgh64HMwUtvwloj0saWnUt+KVVnbWLQhUORLFXkZCLzSIlFSmXMPAR
HUzl2IVqbFhioNrTzzfQpJZxDnAGfHzSlTZ7TcLdwJRHTkFlaYxqQhgN+AlZqhDVSfU2ocFPa3o4
LqZU8wMpEfsWGd8d4IYB9afiE79LPB9tprmQ5v11++FI7ZsfWLouZ01Aw6JxHXOuiQigpmkMUm+Q
0TV9a2wllCo+OEjoj1e0ESYB5VK7HPgTh9LyY1JHPbAeU+E9XPfzklhGM7oOgoHsoagWK1feD+ar
wMOtSKxL3kcNj9pz18VRucptJf7fkrzz4UpX9ZEbWLTtaZDLta35QY1aFYnG333PM4nITbl8WB48
JAmEdQ+IQXY6sRN0djbmH6atXkJasOSiPq+1MTR1FERbgHbRF46IJfgSg4W7ExcIBVZp9HScG5oH
gUy/FRdH+kfx3LKA9qhIsExQpNKj+tzotD5NDGbL3t0wGCYUxeESN7rwwWS4+s2YAoHUzBqlv6R+
K2Q7lFpaGQZsPJst7fgp5jPuiGLheXa9BvMV1d+M8FA4z398eLrLK72ZbrRXMlQtKq3O/05ulq29
jj7q0X/mOzvVZ0hgjub6vLrRtuCeN0fIk4MVUgXHF+x8itMOfQQN2VtgAM22A55rqydmBkDa5MSG
aYTG/jZtZh2RGkZi1hxtA3YWHntmnxUpLclltuy4sngjpZkuezvp8UHvSsme0lVpqcceIWSAp2jw
pAFnxpR38kHrI+3ed6F0MUX0/Oy3o/2h8I5Jlbcvb8jOl0Omm4WWPn3s+lc2CliNtSrgFUZu/wwI
QlKkXX+4Q72IZzfEexFsbq8M8OPgUQAGXC8C7QpDZ+lDSdNIy+5553SV0bSTMNS79ZpVRIPDHmjk
MaJZQnq9Yvk+/6KfLiyYRkJUJUBYtBQDGcSuI7tSRLC9xCMgLGp6DymBrldzfoyFDhZJyd2e8JKo
1YM1M6I9VwC+zC122Nat+bzxNL25bmH7wpcV5viy7m4AZJNWJPmBxQ92bezJfYHcgZOuJyrNdq7F
CZTApCWB0sku3ZwLR52LJvCqrEQv5ZyU3lrrj/o+UJgp49Tv8ZKweTKp1jpYP1in9xyAJFSvlVzH
x4Jxl5KAcGG2+12NpwbYQXJE/CzhhiN19drbobUwQLAvhqK6u4iYab4m+lmP5oTYD4IqnXsQ+Ewj
xkjGoY8mTkCFwLHbs6lI+63bLYtiZwaTD8/OrlXy7+in8LEnzOADuxL9H+FHCCsJyVGLGpq1yl6D
niCopIgT1N+ZJ/pL6IZDf8vilEmLew/+GjJeOoQsENy59z2rynqmj4YUOPZCjJrl5cUYgQRtCMEr
8eMGxD38dzs4VIk77XnlYE7H1H1zhuDXLSA64dC5tXVL86pICHVbeYChUDzLpGE5wI+3F0IgvIIR
lHt3nRbTYsaArkabGBOsrWb3bNnI1jrInyeERbBD+PhQD5/E3cdWa0fpg51w4pPxpzGnstj+BFIR
pQbDzAdmGVk0zT4NFXONvBDp8deqa9f9OSLuPG9+/rSxJ+byeKv9yBVRzS0wl2JpU6NfcN6OC+Wt
ad2uXtw2zSHZW3AVkrbdK0HwGTuUbacfxYz08Ruol4GK/GDFZtmAJcBExqvPsBXxAw/dfkuMOjB5
laOGH5IL96Jc536W13dyDIiLfYKAay2pPHwewohd345BSEQAAKdgEw84kxpLpsrvVurWswXBaORB
LARRIM0a27HJjlGDiGkUaFozu/61TtAbAQ9nT38wPn8hgJGI9ku9xb9keC+99rFVe/ekImzGkfJH
nr5xjtegcA66t7jDDq8PuRBXh8wxenHavE1DF3QgsGH5sSMHDDKuCvPtWYocUMzTsOHWUnEtWWw1
6ono3iUxmQC7PZF7AkVcn/PeNArSQ7a582fSGH6mOMSnYPieNBW8bwcEAAq+HAUzYVANlzGg/jXM
PkqyRaFx7dbLhF/BMQFKafVgMYevcZcSAVN98Le0kes4m6Nne9zRKG8d91M9GLf1Ao3lGF6P/BRI
4pOGIKQsKPB7NjguK/K7CcrvQZ028Hko1J8OPidiXpjreLXFDwG3KT6GxrqTcx9sZzj6xL2F0OWw
19rVf6Y4zqyNU8ve03D7brj8JTjsdIv31jLf1KhmTLY5vjWZsxXNrCA9tZR3+JuWMcZvQXaqkwOs
mHzqRlwyI+URUu7dcgQQxp+6yS5tKDOsd9uBC/sxIGzJ+VIIBogjl5YKyfIHkiOMeQ1GWkxavUtn
nkJ39byuJMXoBZDoXVf/Q4PUzrcm7T21/KAmh/nAhqQVQD3D6e7FNgU9cG8RXE/O27eqX4NcAKrb
zT3kO0EJ/J4pcm/NM7ISnnMXGm5RGCg7A1kcnsI+sJaM3QEuhRofkT3VWcnsMYi4SXT4+ySfKET9
4nJL9x3q3RIKtCVyOSCq+7fq7r0zFZe1243WndeiNKBu2EZayVm71OR/aTYU8FUOMvwe3TC1fDCF
+dLiK4vOm2sTFbisWMiMa7NMZfnnfhyaZsivu9DAkl7HnD4FlnAksNZmbdwAoosknDmpXKutHAcU
6YJmCMUb9e53iCZnaIq622/1ERaKmKpNtkKk9XeXk5vC4/K5/UALqG0N8ZEMPLcwMUmnHRMObyyn
YNQINUeC4tHXX0zUPG73OIaFR2siCd5aC8TKQOd2ZxewTod6CXDwhpvCo90EyZ/RbqkcxeWFOktK
8ULW87hjxy/4mzQEp/eWpd/VjbibEsgTUFWq28VabgLUVAucFfc8+CRnkjeBcCMGT2/Dk76b/Vdz
cNNhOLybqI85shu0wnpbsC4aD5+XLrlfcpdSoGzn3EPgZFrRyAnu6lEklowcbB+5ia5eEM3lIho9
5G3x546DlkUDqk7Nr7plrVu1qZuRu0YFljuudIHMAra4S/bPkj6ZgLRxrJ3Ov/8nKZwazvIpQTtS
TUa++K/rUXfBulPVuL/gGc+s/dvhaEGl6qnecgN1MoFwxUIMzdcsgQhkp44CA7l/uLPr23PAdwsM
MHXFUEmG2aObLshWi8WYrrju2bhTVExdUiTgxWxIqtIAk9vODwfSvnMTu/x24QELFXQc4UanfIwl
ndWhadDNvH3PA3Q7+c/TvUJKtiuodYYAjzNndsR2wEDfh0HgBOG08qsatUGCUN6DM6v6nZbC524g
UZdPlaWydjTpvqxNQizc91kCWNkpqJuffwhXn+nWRi3TrpzTkc0DOPedY+mzEC+O8EtCmW7/H8cG
0uXZYEsmYVAL2m8Zb2yjGtaXteYnCKsiLhso9VPE8gTnua9yJUKJMSZfdDFVRyFgyfAoUeRPrT6v
2Qdz9cOQZvz51DfH0mGLWInLRicp6EgxZ6Qs74+S7H7pp+g584aJDpQwstDxoYbJPoZFcB22eYbc
jPMhD6enpzk81Qpap4UQ/unncib/QHe38FQafsUOzHB/BHALRLmnil+lSAQGS7W/pcpU1xjUZiSn
7u/3Nm0rCmonWGds5Nmsz5w+NL2I21aqe6+VICeJEFevXiikjCu7uKQCFfJv1NtB2Jqn0EOWAkUP
RPl+Yis5eUXaSv+hHa8a+6Af/SWvc4mfVgzJRvKSQZALjxBuHl+4FQKYb9mL6GiXjzHmhs3kLX+x
6MAuQXd1cWpMh8GvF/hC9st97EFoWqSmFHL6YQUmXlDnA96EELesDoi+2YBC/6JsqsN6fxIY+DFS
+WFf0KX8AM84psH42lK063nYtp9X0Sf7Qmf9sh9MzvHFzg5ka1CLc8v8Vson+y+NGamO9eFJwqZ0
ehRxJmRXijvI2kl4JVOObzhsb2tJsTwXsBlPkIxPDJVgh7epD1e4mhozLdmzN6oWIpfyKDWKYZjC
6wsX/CCwg6XVu73nRtoCoyFRJr/c8P+P1CTUAonhb0/OAvoFFA5hboOpKoTygVKMcIL6Bms4VGfj
TtZpIa/js+/PYaggLgpf86GaUqWGkkZ/8vu6J6Os+1CoZzTJ6MxpXW3KN06rPCrOuD6ltUbI4HMw
3Iw8GhZMpUihppAd6o3qatqrYPe/aiCME08s9B006F0Z3XrJzhIG9IXo4Jl//MWFn6TjA8g9345Q
4df0hrOSUPbybMNh771x0s0uHfZ6az2NSu542YQk8h1tyypXnY2XGulM01BpTFkHr2IIhpl6igpd
tJrRINiI5O8bVgTp9msjfmPkm9X5Pdrd8hwsfoBExwNz8vK/CqZvZT5/v7/hEmVe9qfj6HUrVLlp
fdyU2xAdh5ywl6bc6lJZIesKSxatJRx2cd/zC+oLDx+/PdSCcr6dgoktN3iDkSWVteievBtrlHVe
F7HrRmEb9kGITo24kHTDClQ1CxAuiSX3iR5tITp8EMWrZtPMDhs4fa7XtXBZZyXx51Iu5qAiOuN7
dung7VxaG392lziln6JvkVXZdssnAOxVFAlU26vU7sq5RVAgi2l+7No0MN5gWy27CAgJ03oyQdgi
vARb1e0T3wBLnJVPqmWepCIz9XjtAHNNs5JnwO5oxR6jA7QYfsyQVXuMjqo7VampF8iB38K4h+lo
iNonOdYSfovNtfZiJTgAlUCp1E8OVMt53ps2kFy3gMSwgULVHyl2mWVVlf1pFZGLkhtUcee756pp
02FZtUMMz9Z/SItAev2F2gr6dWLl+znNMz5dJ89LySh0WVUw1fgZ31GSxSKCH42sREYSKvotKtTL
78ShlWc7aqguW0OqoQ9AGAvURGAz7a4bqBxlSzi6oCX42TT0sLYWYJ82Uwy3STyXIF3KwMb0qak+
X5q9pUNx3nIv6uFqn1DYAWSDGZcusqeFJ5hRozXETJIWnq+PMbuYHJXbetgK1kJVfZyJLRZpouN2
L4nyVFmr7YSGGA/l4XXhHnhNMkATEOi/q5sxXYL/RefvaE3xKN6lZX3pm6Gcvl+tzQleuRwCrKKt
2ydDwVQrnKgI8ZlkB7jvOXY6DiAhCSIGua+96Rzi1VUU87NryMb9q+f/769CpQcPZJf1btBbxfPI
6ZKuLw/PmQVpDJZYaQP48J/tw1JHNRmdSslk+2QvrqZydSNKVARfRTzekaMr4MQK4rmoSo5BRWR3
4JE+9WTtqffRQ/rYA+BnWvBnKFiM0foNhmBaKW/maWhp2JOKOpVt/gPUZNPZ8xlHk46aJSHabeNl
ki7EoBT6MINApCWHazgEbPwK+LC85kTszjFY6ybUHpfcDjJCAIiiDITzh4AmcuOXGgkLRKsEtdWo
Tz+VAcyR88TroM1rqdU5nFzBHKtlT0uqLyc51835y/aUpWXXaj2Qti0HaFqSlz7ZQILr/Fplak+i
SkQWQrAVPFYeyJ3FZZThn1RlU24IVLDI4x0S/9Da3VqZCX/adZi3su+CCOQtsPTsTmRQvIFP0byz
4xmo63E58wi0NSB27VzfX4D/GaO54F/NkU0ZBrdbWWC1h8OLNEpN90uad0uXTxYPWOLyKwMtX/V1
JBaAbxL0ZeBmBZHUI4FUj2zI23lWnBg+M90h+ifXvmiv3gEyurFCvrl50I7JVRFFYz0uKHetcKff
yb5Mw3IkaWPZTi7w+BZfv7HnInbDMpqCSTs/g/5PB4RlsAK9u7ml84sOIuyt2Ia/+DzlCfTNcwQl
LC03fcplvbLRd7ExyeRtN6JwGWdnKl/eix7i7jsyJeyPQdB0UjNXFBVSj5c8zl5Flx8IBKgdocN4
pScYeAJuBMqnVkQhWNhuVdJeECOm524YJvUUT6RAU68E4IhXvBlxcJ9H9c5s/ObEDvWaHyZ1oiq0
ouDLrr7KYQ+SLJWATrJVo0Ab8hNfwzsforACO4C+1VzObXq2qoT5wUidIxz1pLQGSb9i9tw4OZR2
dv9NOuetbrXnp9W3g8ZvwVvtfM6Oeb8qqfYa+HoA114STv2Am6/uGkFpjfIWpiMHDIuJlYvN4ZUK
L10gs2EcghQnaHkbYejSpBdK3BvIy7qMqxSa2mbOznyFG2TWLeAuoG8YOMkZVhXxc2+HBJ3NOeF1
59UHQC43c+J0ZR82nMqv+FKcoXQKaH1G4jVovRinQqdqDaMXEFRZvPCqMlJqXfHmr0vuvmHkrhPN
nywCVBNR6+PNHQbQOfW8tEeuRb93uuNzla8nzw5XPao9f0CKXK68kqCHziKYboqMflfZu+BMm+jK
bbJnEPm+noMIbgxv2mAXU/Ie5pJKrtjrg3yKnwYD9GBTGCxADHtVFwdB20Nge5rj3bxLG08eEkll
vyjxFS9N6UwQG8D/l6hKsGKR4vOS0IvcvnmV9yiigXKmktKvISB3qHF2+R0evr73lcBjuzwi0XJF
JTRMBjvD5oaHegj2JCu3ovq5MpnZYuE3ePrZtKvExUWytzQoh14fLuAI/9I9Kc3WMH1wFfPkoFHN
4W+vJfQlmxPRX7NYRscdznXralxwrZGqeqxQy0QSPViWBIY49MCAA1wC+9H/lbDCtXRFmwvImosi
bXGgCJCQsxLfLBl5ozs5P+3AfpZZwiOehx6qnGQchOa1v9FhAZRqwk+dCVQ6lwLn9gsqa1ZbfBvJ
XxxjjElI52Fyp/vAoXCXjoZOZdItKTBnXDpRCrdpQ0XT2X5Ju9BKOkNaXpzwRaK6pzVlYBFZSjKr
MnQlMmmy+WIGYggX4Z6THY6nQu1LtxhfF0LysqpHtqLd5cCBNAyTkfQONtmuQPyzy8hM48yI077u
tejK3GJbt5cxZCNziysTFwmoHub8MQrC9KYY5TnpoiTx9v16cDvx+hTRZAQVKSecuduIZiTPlwe9
XYXjHCWh6++1IsL6yE6Eun485fCYzFBUY7+MkvTkPhEEejWtdP7Az405ZjCjEysJDPWXV+JpAGAd
EA1k0+sUtCikIom/HBClaXxrrX/jIeTkGQPOijarpIRmi3WlnhgqyQSUcqyiUjQEU/Tz5MQN4RZF
QKtbv3E5fiYKw7fITis3tc2M4NP3RgC39h8pP55S7zGxjKGpVkU8MRxlDnjtY0mS8inmYpdp4cTX
dy8qNFFK8wdWKeTnNVRl65d+z7dtMGMGqpIH9u7hJjnPm9EGhc5RBo/RE1gxkQDleIvhPxe5U0oo
3mcZKI0lA9QxO7NqRGhjsQi9Mh7MPJmxwRS2B616lkA/qnL7QxSGBLtNzOqY0vh5jyvFks59eYTh
S+49DB5SD9CLQWYz8g+z9ToIFW8BEcmmN9lNkGPR+Hj1M+2NwCaQRwGVSBuuVY5VK0RRsnUSKjzq
/ABadMd+U9RNKz3P4VuwUI9jyYnyrTz35w0TmRy5YrMcfweq7W4jFUgHbXpbrR4RwpKNM5QIhYFo
asX7EbQmZO3hYceWgeBGh5dpa/nvx3FrARqvyfio43xFeH+/zYqmqos7nwo5P/cjhHtgVbEgr/Lg
QPs3U5avTmX46nwrq1wq4N5S1NpdIwslnLKXb49wMkcO4roZXPCIbNft7MIFcFY0QL1PquQ0xUOy
KOgSja5gvsDMYeZNSOj9PYb+PNl2rj10k3LyBaL9YPSd5vlEqm4PW6y12MQsAK+p/syBPG2N99iu
5GNaxvYD/AOQWxcgzdkr6q7cTA6H4bS18rXIG4guQwB2S9XYGPY7lcM06bex1fWyP5bzR/Jsvo70
Zhk1KHLukIh1grf8GO14a39Iod3lDv1Tkl52G0e/ybflbXL5moOglaOYpWsPwNwZkCQK/Z8H7Dyf
TcQgo4s7SUruEVNRfAJ28BDUmGSi579BUBKH07XGStZNfcTJFCt3Mv9rGB8z/mmcl3y4q8Kh1eA8
lTIvUsrXfbNRNLZ5x1OamNdJBCf0LdIb/96znWLVFilCGI8QVk9oSfN4buJk/ILFQUrDTy44ovb7
5/zgAvM/0FcS1+bftmjW74lRu62toQkmjIyPh95OmvD9BbAvipBtuTzPD3bKt7q8LWDWB9Bo6ua0
cBZ0AFlENW3kHf/Gp48fse8xt0//2w36xs+KjXYkxmxnrJOWlTj1YcaIuxtynmQmG5pWk5f5Ry/+
tMXiZdWjPVoXpHXCnlI/Mh0IAjeTgOXd0kUw44fdr7JofRRMzYPURxcBl5S7Bu/zTcE9YR8v1SQi
D15UgnZtnzjndCY3SVWbP7WkYkZ2NMcfBZW5oEyLnovJPKCyGNlLtbemKEDR7y9u35lQE8S7KlNs
f0oJNzpBFCzh67pIHjIG3r+hGeeqriuAFZ21gd5AqvdbFLAayWPhg+ekujMrwD7ts/veLtWjETF8
59g2U37ywfEPBe/IJcMxIRGFI1rA4wMi8FNq+90bhcSkpq7DWKNPhatxxwV593kBIA6SCRwhTtAF
/N6N2bcHbnqYIQgAq15N8DFol8E25Dd03YKIimGMj4p4QFODOqrk9Jtpt2kWlVwVCYvyfpYuDw73
BT3PtvAJN0yN09qCcc7fAY8vlFg3ps7fUoHVyTe6UmonOVKaq0n9S7X1aMfKsA/jiEoUoCi2FFUW
CUFsYTMOfygDjU+pPcULjcclzPxW0mpUxc/YkWGOwmWgOfQcrmYUYwFxG81gH3olfDWFGls4s2wh
46k0NYUHCCcJ29NGwdi0CgtY8O453xYyRe3+1OErzDaSlEEPU3KBui/kk2jd6/hLt368m25DjnRQ
8V4lcZQyN19o4vz+ymfJ92c7KnnSc2f54e6jJ+pohaj4VEF3PaNfO5NieWM2YZRHeQlTWbsqVnFS
tn99yvDRqcXym/8uTXHUFWMVTaBE5R1tNF1MFkXQW11D70DDwr4X9qxSBWfmg/QvU2AGFMbTVMhC
8HOaEv6UgIDrytH9+sKm6DZO+5N43dRnivPOfuc0TUmPzcPkenQFnWKLzDPCcZk6IrJbS7yW/1JX
i5wLe2eP7V0JKV+nL3Dv33HF/CFYNlROnqUajJZ/E5B3Odtb2BjdYCLH9u05kuX0+KxLNJoRCWHH
+anqyOeX58hecSZy9HAa+hjtVuoMH1ZKOO7ogRfkXx62aDlXByCuJn/w5Mhww8AxOPApiYAf1n0a
Sab/YFoMu9xgCdYbSt6NyVO2W0QX2QsZ0DhXeTy5qBjYv0qBy7XEYjhIw7ea3ILO6vTXrtCXfWdw
9IBx4Qyv0i1I6g6kpaNg7TVkdgJCOtIRPSTD3f9IFvw0GAEVTjoinhVKVNVjsb1UBXzJJMjcTr52
tg4WS4WSBNp5NuoqNoUwstqffNvwzii0WJbAbIMXeK4UK9W2016d5dyrICezisZifieCtGVo4XnT
oxZLfc+W2FcbQ0xYwg3xqn4GKlWmRFRGJzFHpz8zXruW4uOMIWboNW33nuW8WkDlBN3mrDvS/t8z
x59IGG0Ur/YuWglESID+dMBkFn0jdyYVpZ5/qbqWrtK8z6rEql3uIG9EIZdrMrCncpqmgkOYxnSB
UTuhs087qjme3z8OxpxTtYr6hQEO+NMWIb1AawibBJ2+6Dd2wp5akhySfHSwTtinNcTlS2NnECWt
88E41gAomxmA0C7w0flQqhu1FE/KyiEkp7U3sYH4dOhi90WghsGfrm75v8kPIg+/o31dcDxI/STZ
fhZ8YWdBA0Y6Y1a+oilFk+Rfpi9p1LcwWz7ZVcKjUMkmcbXdUuaZuWqLqtwJOzUBpUGkCLWvDvuo
/SM8A+yxn5lqdSjg9NH3I75jxh2S0Q7BKB6fxCKs5wSEJkxh8yZEGnckzuLj/6luhMxcW0NRD3Uy
Qj/mBpCAtdrHJDYW9hJpD+/AOsLvYYSjDPgM4LUt2OcNxVCbtDz4XYjwG3vzGHiH1O59grTBYGRe
Lm+swmnTzxE61L+TPmR9d0tFbEk6id9bukTARFBopUC24935hTlH2qeuFLvnCQVLjdYtOkMJj96a
0vQkCaPa3l50IvEx8RscUqfavPTNM8QI39yb+RuSKJ5aR7p94hz0r8+8GhhX4szEW04ZjEDgF+5E
lZJqGYRssSFpPGibSAgbISbpO1y0z00Rnkej37swPWblhrC9us1x2k1oeByg32QYuH8xlVrlhdOG
oyh8i4k8E2jQ6fhgy1gtRZcudD6BwanQd2U71hsnmgY4k4qjSJ3ODZIsXl1MW/xBPo6SmPXjVBYl
LZf9apXJWqFSohfblUqTH95fHa8jD9IaqfWC5T2H5L7eLyVDo/WUogpHYyTOAlSYRNRJ9gpIBrAM
qmX01XqqF4t3h31MUG/UATA6e6xpLM9Mt1HFqBy6bdj2fDWVPc90INxFv9VdYsLKOWxD4FzadaEG
rSREwkM0pOc6NHkC4/lUbhIejCgxpXlc/jGwkIkwoUH7vaKSIK5o0gWEssuZZzEiRjTRnT25RHeJ
F7G1ZUj6a5WNe86rOj1T3t6bBNsobHK8TvCrdpxLTEOErL1L+E0crwO00YOOd+5LBW1jp2wNGZ3l
JK0ZtDLHLLGTxqHdNwEoT6pXn2poK4oRhM8waj33RkJIpd+sEwaS5jEKSgg7rrW2+FQgff78K2Sj
wPQdm3eH67x4LR0emdO0VoKrXPMeD/xxu8YMJ/f/XgHhM4nvzIaJ/cRisQwk01mRfSATzvv20HQm
F33eeqrawXgB3EPYfvSdSfAy4lz/A28PCxPjWE7mk77Xz0Z6oNs00KljNuXkGU92HdQQGyb5MHBh
FonKYQu02UMotih5yjT9BMChCmFcNV9mAeqWg8Wfk2/zJmRK8wkOEZu1a5NnLKJE74T6F97oWyyz
Di5VF74BfLdr6LgqVLMmcfvWQ0EUJdEfS2KQmfY9zbBtyooUUpbUQaaaqGkK11yTLmH8pZDQKp6N
lWXk8ckcTgedd0xesTPL2MCKSZK5nIIVuNHnAFhCIquHFJW5jPLV6CStuGK8Bd0g8sVVLzoL/lei
WI9dIs7qLzENpf37w7JuEQyxhb0lGgScfh2hZcF318/I9h2hqSjKYyS26BkYKP9hFey2PZKH7lHH
MJgYSqhBuvwVmkuecPwoDfTSoBVHuc9n1iKAPGCiD8dNu3TQkbedscE/4JJRC6WtNRRwMIRV2Svv
5cLKh80P9ZOYnzRhZfvwQdDVXgTO7Gsp7mXk/1HfG1lqempSSnUMjS7r4GKiB3Br+nVbulAT1Qal
I/x93Wx2AYqZl2lC0cDztqG9nWzWrWpkqa12C40M+NlCfbpSxmGGtmTyENF5JoYfdJg2xafMDDmO
4B1dJgsUg0K5/KjIChAi7B81Ru3YHvH9ZBXptdCrQqitJndlG3HsQlzgTDxwlJFJUznitrqjDUTt
eGNwl3JHtuqX5ZCIfRt6V1pfBeAxfr0VImb6v94pJn7xProrHKT/ZWWs5Y67yJYL3gKNwSUQqVdb
SGY1Og96zIi4KOE0gRFUNjHuWDHp5pO5wL5Oyjb9ej0T7Zzmafbs5Dn9JwxIW36tF3u4UdKUnVgf
hF6+L1DbGBZt0d8bQnec1EWH3JclesiMykJi2VB1Df+bfjLiEHkUZ3W05PVuGUkCAqcSeRPuHdmv
MLrT7dP6BUBjKJ0YoVxXLoC0ZtGSiycYug89RYlcpSJ+2jbOZnoFUK0KL6NMNISpuAib0zU6hTOT
H4UXnhLXqbCEp+Wm3E29WK/Ccesv7+4o4j0EJYcnPPC8n0qBufTtTZrvWZn0nwoFVQlabrYLD/VO
Hf4mmIBUUW7/3f+7D5gGMFi6xXL7cSln+wSdTF8leOEEyRAuugBOt4FkBMLsu1J0PCwPnPSXJKgU
zr45djPfZ/TZCU02yd3ZehlWMvvS1slmPbxciH8gzU3BaeJGUDHZaJ6uJnYnDVl+g9pJIAb6lhJe
yrwPk7/7hWQv/2aMMkj/JFNtiCGyib+F7GD2gncatwxDQaWdypNIGyWFtFRlv6B67qnVO/g45U2J
f2Uq3Kn44yI9lXLSwRpXRa0C3FfwGnnR+quWlM7UIND3cv5EebvZJh5kTmauZiVwuWGz2l+v2v3+
Wvmri7ad/AMjtOya87sJDwNVi9UJoxhs2iJ3VQJrNRjTn7jQxZLZxxoTbb/DWeMMKneGktFml9zd
GTEZ0U5POqhE6k3MTu0G7H8xmHAXG9abABE7A6mbvRo+dfQ8sIHMXjV9Tun7pSJwYmvfSd1OvoU+
HdT8fOkLrZ8DA5e9v4+320SdG/Z4miCtJzLuk7YK4pJiTiZp3oDU920ekVymBIIfoNxqylNTOcpa
8cYvY4SgQ2NHFKe5c6kwtAOtB/9ZrFAl7J+NLoWAvF7x4oZ62+R/r5E4psGEMKjn6+wxdfBPZQJp
PwU2Aif9bFRCvSVgH9HCpS0LevgdA15EjlCzobviPjswFE3WWP9+1ZWCzn2gMG6HxZJyZ7K0uJKd
dw+MMhnNWUwy6Ftx9P+L/wUxSggEFaMTGgBdmS6mFuAeCYQuSzkmtN1wMOawytROcbdV/JpKhJeQ
msONjemRI0y0q8JanwM8YMEQXNMwr5OBqxY5tKKfnj0WlHXjZrCr6WbXBxUdAZj7+0kp7qxxnfMu
Ys6V0cq2mpC4fJqkBR46lOPbweavmKMd85Dw2WDBEQ34A2ANXOCpfBwqNItCSJX2IFn/4DPIwpGL
S0eo+Q0HBXpqMDM/hDexfPTjisxat0VuK8KAx/JrEIgdSNS62U+AhOGWMYj197478UQG+YxT2knm
CzvSumoXNuu+zQLdGcXJgeqcdtegirgCmJ7MtlkIIVjhjGWHOwp0/pJVHKRM1qQaCvjH63fhnE3q
/ai4QIae6DO01mG9DGuyk9XBSlXBwnRKlIxMtFvbj932oUCvVOLdrDWM8g5WKvwsql8YnuAfPtgy
e1ua6QMn6gF4nf3mGN17cSgCiANFDxZMEBzj/O/6zW3fnN/RKD+3an1IkqRJHBtcqi/zIcpWSXvb
yZz+iJRx325kCGoUM0kqOvGEPVUrAri48nG/Df7O5+iOyz8u5mgqGQ000s432WurlTswTTIwlNdK
IZ9FUmizliqIc4QJ7k4jPvDeKxzMEb19LnxqNm45UpVdvedrWBiw5ejdYP5jxKw0ZaWHuHvbeU1T
mhaYvrKOEXVOyj5yy9D7/StkkcGfCZpXar7Bah/TsrWNEMG8gzJGUX53IZiGb0UV89vSrfBuvL9b
6+vP7nhDw17wlfGQaknWtJOYY4HGzjAxWsJZvMoKgOQf0NTp/BI9I1GuJ/T2syCNhVOGt78vEjYF
C4KmuDNV/pZVV1E/y5jc9+KwFiaUGLkLLhSzAWQ2Z+NVU7fccJpoXz0vOswIzFyDDmNTcb9sbHSM
/Kw16XEFqKn/7mCGgcoqoOVwoDYs6zWa8sG5Wx0ENokO8HAofLiAf7ac2duSGK0qBBONhv37/CAf
qv1QffEpkb/TIQooz5x5iohkUE5CgKu4/1B648PmZqR6pHidZjq5/+NkHQH8TO2Hf4VT7g4WAURy
/vw+76J9Npb8gic/gAYK8L7qy9/z+mWvw8j/GqZ3qa/auWQDwTJK9kvWZVP0BiOBhkazCl/DB5Zp
At8olPr/QPPrEZybA887pautkMDVSgDOqLg1WFvUNAu/FFvcReMcBIpqHkEXgrBln0z8UgzQpDpA
1WJxxfy+wg8KXI9FFbaQ4Guf+UFnBTLUBJONpRRrjAgWPCUdKGLYuF7VUGkETb9g2z6bmvktsNET
ruyyKc9OgHWE4L4IS2KmmMOsLUcpqIoU/NRgLAYezFxJcVhmXX7kCWfJTYy4duWRIBr6a2kZgQMk
zmvhgRSAUU8exTGKWnT7vWCPcBr8AYp5zjSOdHhEUhWq5EJzyyeYX0+a/RI49+5d90bHZj/I32oF
ZXKRB96nLN6E/YWSfzRC9n0OTwL6cbpaJFnxMpiwzKzuKAsdpMTs/G2pij6c4ogmeLCKumJ4H3Sr
pUbC7zFFAVK3dck5zNs2nAfZYzuO60gbB3DTlhTjymTaCLv+5Z8xEj7v4LNdSukQKt6fcXCNZrLv
q0Lls+E8H3Bycw0a2LdyPa5BVxMzFUIVJVNPWfFRlpOvttiPzkkqS0xYsnuOchhnOx3qSa1b8+mM
ml6u/5mZlWEUCPEKBUj7VC5INaJUZHCVzDXm9OZ7+LoDDTyu/ghY8cy78QKCpYvlRmiHn0cSj4XK
HDXNZN9TFEb73+1IRa4FC0OaMmKuq6BOIQF5UE/AVJJ2kzQPQQdhnolbqkuGP27DT7dTvIYBuVKr
oj4rqMbCivQjjYE+Rs5g+P6tYr5RZ1AxZtaIoTc+iqLIseTHRBCjYYKtxDBjgzLj3EL9NWVMQtjZ
/YBLRG//EGAP6eRIVvAh8hPgGEUmyIt06ETIDdOebMY7mwBfSB3jhNK/OMvnu66PfEAFrqvhpvE4
Iw6+aJxhDlQyU5m/Tt34uDgAH0vG6hn8tGDnoEGcKuQbMBTyjbSTBiai6EpKEh6tpd0y/cjVCe0r
XyYmY2hVh6HPgv/s1+59l0WxcSmKY5NBVyhxT5DmUJUwXswjafb167/UpjO2nEfUSDXPgleHgqh3
+spqkYT7E4C4JQM8upzpgBJI93yJ3/QKAkDt5awxFF7F4mAL1E3NzTBL+Q44DuMHWB0fxs83X1t3
yPkTX66GqxLQpbw5oEkCNw04nP7zxZgSf5MvBwF7FrFNphvfA9V+/LABWIhiFPU8iJbVHl8z7Ttl
WJZ1SFSVng38pBcxqSolNQOtl1ioa0KEOd8/p7ZaCDuW5kCPFiFQaM5ZdDV3pqCRF23OF7BnHW8l
2bUa4vzO/IXzBHR4WQnILkpytqec+B8iGSVIuifflcd1N3y4NtC0vcKFfMeFQkieq0p4fGMNp+pL
QojrI7PuaCyZ0+zL7ZgHEl3KJEZaZvN6reNVwYAd+mtCHoT1veKJ93xiLiaCE1u5v1rwCAUGYgXq
jPuRLWfhIbpW6AFDEBybulrj6qCDxYy/5L2KUNWjuSQ24287kpJtWMUZ5DSZbX5mAxHhU90gAD5W
xHog98xosX6m/zXPikW72s4vSPARFTl8gihIMVrHwiaZypzykmcF7vfJYrV+j9NBov1KADGqWb+y
Vw0/l+2rlSlDptDbVJdjaXHx9ACF7beFsxG5EZg1Mn5jv37yhGjm3Mui7IhxB2eqM8hZCfVFOV00
ohmwiuhkQjA2Xr84eHvNKpCu3Rg/rC2g4q1HZfaxYDzCSvqejOOwUuCljSpAC3Mu4R7sRU3lhrxe
C/JAQmgvWbQaEqzznbSFLzYsDjj7LOilx8l5DpOLN1g9kex2kpQDDYPkQbitQ4iyI0MBad20EoKI
94epvLLhx/XYoq+gR7tAIEk4ecEP3MU3yUc2mvMEifABETXSgkBI9jXAwEVtVcwxNfLzMmyUuB3e
A4nzP9ceo9Pdb8vc8Zwi7NqcHaDQlj65VGPt3pttCHq3LJnaMdGXVhyF3WFxeR+J6FM9+YAT5cZq
AxJglEFE+o2KRICOn/AwQoo7tuTg8lveaZQF3Xh6veIleBqO2qD4vujkvpGSWvpAjgw6MbQPa606
qZ+ZYFx2G14AbLQIwEEvPokho1G4w127rnfGNslQ4v1Jinq1BMsNvcvu88o1rNIpz3C5s13BldAn
w/rXizcyV6ZsTnc0PXz3vbrfsJOsTYeViy3DlTHQSHaFrcUnsUqmV93L5t9pQUXAlkijvA79Vf4U
9g16eUQFXCILQtMBV1ktfaczj55IoqxK//7qQCO/9cJMkgc22ze4GHKCK0BHbPpy6LmlNYOymW12
HgIwPi7Ln+KQkNp4gmRBdp+kPOyzM4y5eV4TORlCZykQvdqWvPiQ2zz2B1upe5SV8X5rQNp36y9i
Uc+ZGbv2kcwulWIHCRN5gLd3BFv7KzHQp1EIl2PRr8s+QRkUBZMOb4vLkusBBDkK0In0T01NQxkN
/ud1+g444XSgd4FgrIIkvqNjOVtlxBgXw2DGo6BH/wQ/VLH6VbkDc+6hBW3aRh5rsYRq3NrTDs5u
vbPj3wiozbQBAz1ufmI60bJhPxSFSjC27uwNAmYAspfzkE1DClHIKthD+Le0NrK5ryczHQ9X0SvH
xUW7QdO6QeRcnrNEd7Zirr5oX2sJ2fCdnXtccUkyx26UzEFtk99PLsD9MhGoaYC9bf4b0/b7lApw
wpucWY1K75d24I9+sYlqaI6JoZUQoO5Q+AcmU2qQJGir97FNjAXCFY4dJ3RrtqGrY/f6nIjfCkXS
myECYzEVYKr+w3c6T6awZMvvpbpwz/gFWOEey3bJtkxOS6tEdocyNAOr8S7VIHAzV0ocrJqUIY+p
udEPP/fp5bIC9+jdbYRPjVmr9BAqOR5wv0TYOssmoxl3GOQrHHkv/HsOTBhR3aiz1b8Q0QSLzx+n
i641WwCyQASn5OfSavc8bN5VelujRZX1vSItP0/9uJ3tu9SrBP0OiKfa5ZjlvlJ26auHPmOJSGN3
Iyx42RzoH8Se/D9Zz/5ebBlhQV1iDHsiumS2haSO2/4rug7oBfdW0Ko4t52VfFLpH3XnNOV5wIlE
sGmWddhp5LIKgO+7MgxR9cF+6LkdD53jN+GwZC4H0O1cvFM5tYatiFllXSEmnZbR6U5POM2/GnOy
m1FfQTk9uGheI2/OCRSqQrDBt06+k4UXPgsvv4LY0XFi8uhljwCVixwrK4B15GgN64cW2nIhxUZF
weG0XqxCz5+GqvMMZh4loVYKOSrsEqFz/S2y+cz5nguYrWjo/CS0QlLG7iEhWQbWtnuNUkReEI8X
uGB4fLVw0cbbLS8pviINYvkYSW0AcL9UiAGiulAzvakvjlKVUEk0NccQlZnM6RQuxTMcR/yU3qmI
o8XBzUpsgcFeVLhvClVCje1mhig722r7wyioiebkatVyOySQuVft9gNsKX8/KaD+kGFM1FvCJd9J
2DmNqaeqGkNJixJD1bQvVmlAgu3cru/+TkFXAYQNNQOkU0KXiC0ylP4V+fME96TCVGjgYlol2Pok
l4g5E4ASoOZDkb4rTKMmfI6nbtxipW0PYSS8VqiU7PdmgVPzjYkZhR8ukP0C7VOo/LE1jmuviazr
TnzPEB9cTOBUvjGRmif2KKtbI+GwYRu7h7WbcRXSkZGtN7HHF7KIyRh5cR/rAFRQRHcdTdPBfbwt
xhQ69fqnukrhPfpCAr+36EbgVrx7NuxX7EbE7vkFAAcN4huY+BDc3ksv8K72fFSnPzn3nVIWpp+i
ZSa8ICOjJjvACX9F7yncVJfq3WupCGUaEdATpqUBiJyi2ADAWVWjAJF8xI46SE2dN63HDwxl2r5i
8hTuIUXxKWpCs3cLY8mKAwRkidzgTq30mVKjZTX1iHHj7Ci0KMkJgY3QpFvD2l1IGUmxrsHhz+mY
xOB5uO+bJqgIjT+doxdqRCtdY9eBODEQKtsh/oTQ2+olIwZyZ5fBdjdwXU0KTY+YggjXf6/AoQ2b
bnC29H18d9IV14tc6jugD4FfwqLkmKo/Y9MbrkJNhQWP/Z63xeqy3i/p9cazf05LlqztIkeF+dba
1FHdZWRGrM7bFQXnIzibRd16VUr7L0312B3PKMfDnQdznj/k4WCDq//uoFGnCSabF7k6F8B6217I
JdOqdBlQxCoWRT3uqASRcSkDnAb95EDQm+qsR4xZr4cP9NUO5tBb0W0r7EK5MpT9DDY7yiy4mVd9
1RF1SI7d5fF3dhlAZVmag4F4XUboIN9J5ZYmTuCEjx7SXXaAMfB3YiUGoK5jG5nINf1nJGABYvp6
bMVjEDSzFlosjyGXkmITtdZQoWe6jFlvhgNnqnVfpw4Twnm1+VHCobpeRdp1VjcbBkS4ivr8Rc44
Cn5x3FUee3tiHKoWCtc1ZwMe1qJjM2/RMdD3C0WlkozjUK+wrCx7LHEPawf13pcMntE8VJ5xcb+z
UR7+hCwat3WO7OocFnHJW05TYYS0AklbagAS/PLgKkAiGSrDpYT7m0wdcnzK7mQ1dCIOz5CX/TW0
2WRo8Sck/HJIxMtzRlX8NnBhs7UNoJmjBkeNo5omZGtpzHqOLpzx26lbBx3CiCU/Cssh776YXQZh
BNkFrrSJSzzbbW+ibGsdJlN78PUA0L0Ro5gbVzXXT+WJvTjlpqm4/gwMt2xSkk5WKBO6ZZCQ301m
R8f/u1546DY675YS/uLK2kdD3NnNLkc7YywmNNau3jvbSmhMae05RrmqbJMjdJ54j8zss+vttWMx
Ni4Pvsg0DXoT8+WBE9h5yIGed3k9tBnVADzzUUQiGFnEVXAWk/2FXrKMiXC6n2QcOIfcMfevQNII
YYBd+8osrtKP02ElpwU01fVO2S/VlE7aZ4/vcUS6QD8sqE7ziS7CUFpV2DmPWrrW5MpLa0zJdNIE
a6oFrODH3RHUmNwc+iptwNvkw9OhWgQrPcKTiyvtvYwgZeN6DQt3Tj0ER+leIFCGKCM9/sMv8e7s
6WMa0hWgl1wIIziyAM/Uaey0Y24ef5L5JetTALH5jm0qs26FavhY9bgXKwGysZH3OrKJVJWN9jsK
7GRQN2SdN+i53UUtcDYijjn1/O6/zCIQd/yzxOkLpynoO1UaN+cW6sXjS727ajlBBCZt4/7g3WQ7
P5+xyiotEmhHVbOQ7PdgmIlCZUQ2cfopYqFpeLTxCAv1gM7gQN3tPLVz+veNXCQF8zlVa6JV+5lG
DaSXln8L9iwoGmmVZzc2hG2H3HAOIrmJ4m8o9wnYvB+Rbr1tVvzGqT8oqBrzbOj4VtuzGIGBxMQS
7hQZUlSF+NgwFdFlhXTOiQBhpiOKq+d/Y+d3N0hzmuYElXuD2aEb1A3YI8qRxxf4W44DzUX7FfN1
I861o3AFXLMQXJzqckVI3la8Z1j5YanVvQRYim15KGEaYi77A2rh4a/4/siPvbQ0IYWGC9gAXVIQ
QXtGIom4bGZlecQVvpOtRjkjIkiSv8Gg69P+71XF23U2Il/V3tkRyZWdElWpDufDVS8ChCwKPWW2
5FTNvzCm2l9ZNdaLbr8MLOlBas4KtpbhSWPs2cAXQ/eXIP2k6jqj1dmCqXz4ttrV7n2Nw4y4l+iz
Ct7u6RZq2mvOSI0LrxP2yABqv9v3ubkZHiif5muflOK+RtGMMHO6E7M2P9LUdIRteJEhaXFQ4NyZ
qOGUfgVdHLpss3RYvxmZ1lPlEzRKXqKYbsYmxc/vGca8d+y/nOWyLrrDoIWt89LEFY9XxJ4cOHFh
5bKWMDZSV4/90/MyZiUjgcBxFPBqdpmrK1lUvpdcGbg0uU+COan7WvFWy2934itR5yzgocc+3hV1
xUOg0K03vVT+GDk8/hEbkix11UdSCWk1iSGQkDEjnjScGeBc7nRvlLZgR+5Gy3nDNll9HQRgKyau
wADgyKiL0w5t4rZ6Zp0Nixtu8UoiYeErBC1jOn1E9Od4se9BnFNI4lZTNY/7VRaCzAuSIl+Y2JAo
Fb4AL+kGLejLn87ua8d2RECIgYVv8ceW7sPNZwUyUiBdIv55d6rZtWu5qvpDwbmui7RnXyXtt90g
ZNaWb9KEBW1tpbQhn0Ti1XuBJTEGx+GammessUJcLz1L+9JgNoZn4XEkCs6pHTG6n66sO+40HpdC
ZOX4uC+1zfV6L16FKPtLmVG7DuR5KK1IpGcOkRK3ae+b0yQFRfwTLWgNC72gkmbw6kTED+t+JRS/
RWL0Ndfz2o9CJ5xZLZeQUZM5k17a+yiqBokqFsQu9WgM1asWtGdBN/pnh1TpLDIFW7PNmYvDupXt
qNu35t8IihAgEqDaL6LQ+EX5nGzfCkzad91qnjoZuxIRSz9lQT0QqEoVi4hSW3VhHuMl3ECiGw6C
7X3K95lT30ly6Y+rti1pMWb9skwQblLE9hh358e7f8X4OgzPz1IZlcFBDrD09Y6PNF+CXzk87yWI
DylKmqSBvcDwHKUep7iOwQByhRKWIOC6b7eFkmXPtHZ8mn7D2glHTXkBANDK2QNBxK6rGqxEi3Uo
aC1B8BFAEK3g/X9KUARgs9GSW1X35+EUFnNsvPcvU8gt8fJEAmjpEFwKjWw9VgNyThl8M+3BuZUb
J2SC1FgMcDDaVyr0diWvr+gy0ynIAkIuETw/5sMa5NiXFFWrGTbG95slY4v/51lAm36S2vA1ZRTh
eIUavcWyg+AT2OzyDoLsQMDF6ebobApGzJQxjBZzJ352QCV3OI6LQxCyWR4PuPT/Yi/vYYvJXvEa
tFUMCD9URbtXFZDJGg9RseY+FxHqmfC5ykBWKomcdyh3JIUz55Gf1cz5CUuVUfX3mNZqzUzKweO0
F2qBOfjwStX7ylPV5tc0XKFCLj6matXoQbrGl351DgalgPLE4rp8Xj7FcuHkDWcD5Y254w2ajS0s
XdCp83Vpp2eqh7dGV2HLSrPcsUIV5Syf7EO8YCJe/OHmDlx8swquA3vcCAw7NZGOrbLcu+bfE0EG
NqocJJVgywVmeXxS7wcshAodvwa+aM4YN31pJced3FPySWE1gCLD8PkBPXhxE8ZjpCLFtQ5sGvh3
GarpwD8gAWKjdmongfWsVDeza8NkUJRWAUnKj/xir3LaOdQcHka7l2770HGbcuEHyS+hTiBRJnKi
QuIVo8uAfkDUEK2BkMyhZJ8GZDGVGaweiLK/JGZ9pQIpdv5Zzwi1/26ATYhIn6VO+MUcyVzuO+nX
m45Hv5RwURZvm0SuNgF6SpgRseRnT1eAXPe6E0fyM+dJhcdesggq2cDG4knRYXwuIcGd/Hl2Vl/O
y2NFrOHOdShTvEVVaUawvPZwnYwM8Rd6EA/jhlR107wxHUJUtUYz5bj9CGUkZDDjHoSWvVHVkbnH
rrSTvQ43QF273os90tSeA16kOivO22P7bXzjBx5TMsRamQw3FvQtNI0MCJ0gJyepW6rqmz38Fvdn
7O/YchyvYYE5EHSvzNFnbKJVbasf/UCPLvhRW8hXJwQe/IXlLO21+VFkRXzzOix1gd0adWtxVeB2
rMgd4eO81PNk2PwyyeM+CK2GGJXlqjb18IRXkJkVYh98Ho85PMx7J4wKOiNJKP7DnNGEI1fib5PD
XZkCR7/3dj867TTLe02z4NrHZFceWHi7C7B8pjZQSnI0KdBVrwz0Xf2z1C6o0H4PRpboOB2uoSys
GN8tWFAgBGp7OUOEkDI/9cZ1H74JbIp0CP1Z0pKmfRWLIKgY8cxkC1q0+YVvwFl6O//0VMfTURLR
xI8JkOyPEyjQE1hPldnEi3bqmfT/CHDJRdpkBIIg54ovEwyK6xhYQMecW0II2d0W72AI/jLS9+IO
zD+tcF4mAhsVoiS5nvChPBtmxB2pN/g0gUTdsgy5VX5E4sNtBn0dNCKSbGs1NECfQ28M4HL5myC0
W4iZXUPUmj9o41wxHhU3YG5plZib7GoLzgAg/6f3O+ulKkqPqRjr6XnOTLWaakeLQlhMSCoC4VwA
pFw/0lXTfuzny4kWhkJrKPPJgPfuyXMz4wX3fGUQa36Fc21eisE3qOQrWBa5Lh8Vvq9lXR+p//qu
bWRV/dJ7TX9ekp/BsNIPI9mOdgOglsX+1E4K6MySSJ9kD8W4HGECXkRHo8Jn5sILAtUts7gjo5d+
+3O9LUpLgNCZE/uJgWNpCfXthZBl/wk8t6k5YoupAINnRaByZcOp8ITdSb/gtQuH3YYB1h16JwC/
YS+Ptp2pX8fPcqckzOvuqe59OhpmNYJKDuWqZNlXg7wDTOOAFj2gaDu2N18llCX9WZ+nLBVCjjjp
Chq/YYAAqUDTjoxPt42qfXoXvlBORqwF4zOmd02Ug4Fd4ZY/rFBYqj80rLlNZvH5Kl0zI3psniBX
hJeel3psb/jFKOKb7MR2Ahpcyf7KWLYXhcDsltKjKey5o8KTC1pyNuU0UfbrYJShfu4gX8wLTCG+
K2v7mI4qO3QRyyoOY3Tg9AMZvyvvZB2W6n9pCr9nWzDJc/ysuZAM83yT6cEK/bL4wcdZTmkD58oc
gQjFVRQXwzoetRkQYcIssJYf6tq23Y/3TAsVmYFYIl3+zCGSSLBKdg3oPgaFAlDcZE4AXrJFquZA
gNz/TEIK1iBMKQa9uha66BGM/c7fRmcEEuv5JBgU404Cra8tWGAt052JhgRXlosylbuA7tCpQyBm
efPAalwV/cdr7QAusMgZ5o/oX9u7diTTL2pI8Cas2LyeuC4lh9Ds+KLN7YYwW63kZ4Ig4YDp5drg
H2bRoEK7OraXAytaOtSedP0pc2zOBhYiG7SJSIRqbjnZvbRqU7En0JqjIFtX8JsHP8IEIKCAz/MG
ZIl3AsVFZAkfOXUXmc+glS1wj8Sv/8EPi+YzApynpnahbYnc0J8+7yZ3rwhW/39y5H9mEQP4uFur
TBCnXK+2Lr3lFh/IcScjo10No1vjq1lbfAhlxqDEwjGZWm/NHM04yg5tyb22ZqlPKGsMnBRxDibP
Zs527+UcnSmJhWSDhmwL9AceI54VHBicxkJFE1wt95jo4YbF34yv9U8a/S0eVCWwamugIM5x4EJb
QnGONgUln4Wggd6WJWyDf6XYUFnMldZ1o1+98iXteJZRozORGEnAim/FCfO+WDTzDB7urtnhOViQ
xM1oqwkbZQtHGCUQHAOGdGlsOIZL0Jmtx2rRRezfMYhaeQFunjP+iItZwyZ7KR1Sy/Bvk3DrAkG8
KJr9WHdP7mQ6T6lBfSSW1jsNEC0vQ7mMWT6J0m4t6ZytQZvdgRStOGkZcfmbaNesomsxECvjeQso
qRmH8nFTNzg0cQLjHyZEqh7E6/37Gsf7HPcQ8SCziHn4sCmKXcIrZHcZ9sq+SFYo5X749DePyq6S
uO8limZX5skTtOgbD2T7y/PW/UJWIa1HuQ6NQ6o5b46N3KZHVEpf9mHI1yqwqQE3UcJ4dCFJrgj7
7qKSoPmsO0ZkWzBUr84voDMJAMnzYHyBtSD5GVAx+hqy4JoTa2NhV/zHab8FKvQnhZq18FoMXN9e
TvXqmrkTTyYhy8lIXLQufUxP24DqtDO9fU4DdTpcTx7m0GQR8ch39xQHObRUrdnAazEJnpbDnvHP
nOCRFZFZl3yJg00wFwUXONqgf/Bdd7+szGk5324EuwUiFZhNaWXEfPfeO/fhaeCsm77bJJ+HrIyI
ZIrLSQoiX6gNJIPJ5f4NBfMS15GFSIR1kjh9mvduPGQ17k3j2hrfPoa1VWAGLDW78nxyRb36EtQl
Wj2ZLwCZaeTdyA2C4UUFgioyG5aG40TgtKuWi5i/Z2WZdmhPx8ZW+4vCfeyz6QQ/RipT7I4ehfFU
aP3r2rZ437wX28uZfOlreXpc0D0em+wxPh2KH6w2qG0OFSl1pVccLOchH5adDPRpfr0carelxRok
AekRIGwXXfk+hR0cW74/q+9rJAAYpMHod7b+6imGNgARkMpZKxdHU/D60m96AdlwV6jWjp8eHzkU
a/99KVRp3Npzc7qPUkgFnPZWhc0ARveycRzqz19mhghXnytiOjGzGlwttG+ULLlgMvT/hnlmmpI8
5CnoMncSgJRhGRUsu7dxHAEMUCAHN5t1MJ+s5vfcF6uGmi+Fum2TGp8ByEw4IgtyJaPcHNbUgK4x
3j01rRRh21Sc4Kw/Z3XWfbDNz2DkwEFiZQuI8a2H2Jwl9/n74ENY8TMC7XxjMB4GR9vExdQwVREJ
agDC2ako9wY3otck48WzSu72ZPHK2C7fi3dxxqbtmER2WABcfHfMarkpVyuEa0lKGmu2Yr2pDHE1
rFdToR3tddq0IFxxxTybff8COQKvbB/gjRn5S2PrOgKI9yJqAP99OS4GsKADaUxyqKwZVvwNqtkw
nPl8TU63GWhQPouSJ4O3hWdrqGfhcYtl/YBZ06QHExQrjXr97tW1DhWXK1QLMn3bHA7+MU44Oht1
TMZaoL5x6sqq15C2u8qFVNPWlx5lwCoXhm13NEdjz6FgnAXIIzuOnHnxUKGR3PArh6O6T9+fPTua
yNy8q0dYdR6gwIqoPaZslmKYZO2XmuQM8aI2om+t7GLCVTP1ImowDZ01PQ6P+1Ys49pjSHIaJudx
vnsP/XFJR/VC/9oQgrxWFpeAqVudsFFxr8m01u6kbLBfoVOBsRtUIDGaOwW4jBOIBN0Jz3GNxL0W
UUiGR8iNaNkalpZZYk8c7tHS/tKnV+6yReFqJp8fCIF6lT67YlIsb7wOKc3J8hdynREJWlI7+1Nw
7xAfwvIWqyuL8tdzBX3e2X2F1QYQGjCTT4pxzl4HN3mRfc/7JhyKvLNmJ0I2uNzNWzaLIPfagqH8
yHvjPVAztuCoNvfJTAjc1j6mfnjFItHjY22spf8bqNK6NjKGk7PCPybLLtCeZPcQwnKYMr9cDAAN
sEshD19I1G8xOg8zHNbtX6FPsvcWY77gdkHMNpCOMKoHfmjhxBDPyhNZ9c4hodcQWn1j+UrtWRvl
1UIaYRmvcC9Irzy3WFQGPDU3nmGTVIRBQr521lrDHxpflPUuxJkMJKBM4uuddraihVu8G8yqclOs
un281SaGLz2ZctQm5JpV2JdkgnhUgHHoFAlvBGu8HLaUUOzK92gFTVJUiEmm6h5vDVTFv0Mjc7rL
y4yN4DawL8kPFLjXBHOzU7CcrpflcSkiWDiecZIoZYonFrMob9eRzcC56s8gvjslJMTwRHwkjm32
v8sp6fDeyMNkqRbxTOYjDqVS9dBOX6M5qqXVHB7ZyVLk53Iqi4YMbE/gBWlzOcSE36h7fTElFuIW
VH2/faUt0IG3LhRu9Dbq4rAomfIn83PZf//Lt9ybK3dFtBMw0LOmvpOpo4AZFREER3AmtvKGWySx
VsaOthxOgIAHfApLVMhyw9UYxJZDo+txtFQOEoHipJvCb3EcwDdODB3ug4Ts74u8A1PdCmCivpwT
9Uvzgj/+ldnl+XpvpGAYBV/8CreYsG8tEHCMd9SOfdh2vD7UUHW4U9NXHcM/hOWYPpwdkkLQgGX7
as1ejzvrjBZtS6nmkJuwqLFvT5BiTh6W70GxSz5JRwMBigU1anmIsYJQgB12DHche+4rKXlgmzSg
sGetm6ypS84UqZ4Cwib6bDupM4+0PFLm5xkibLvnlQjieQmSxHcLCUE3y7zmXTRulWEFKRlZuN6g
3LG5xxMTjhPeh6WQne/wgzIQM04fOKUNeG1QoiJDPp/nl+NqhR9EKEjyS4lmbt2QyC40tNSGL0Nv
iLCQv2q7m3kdYYK57F5rrjduyszVFY26zHaMhXmaXWajw87Wbq/1QjxB8E9qojTS3DbsbnRVn9b4
v1gS7nWeHVh21yhqc71mvDXEHbnx1AGJLuS7zDpDQ0ZE2tBiAaXqFeSlzx6tsSFfT6USSf/dZ1GE
Irtv4FG7XvTfYUKONTlpu6dV8FAK90FBaAq9i0gR7iZuGexnMy+3N08n8GrF8oDKz7i44I+EiBh+
wYHS5SIjnQfwMXqG4GjB7SYv1osNDw4vjJYLZi9wpk0xCg98byQrmT623U8oJxoZvqXLElNAYYDi
nqIzPiw6YF3UxJn5kILbAtnW8aSEwNYO8javl41QjoeY0QIXFf3MyXMuB8urrJcoE495XAHVZf6u
pbuauk86YNywJX5wcepw/Yw2zQTyi6D7ISpYR0SSd3HP/TIWclKfSztP0N9vDo11laB+htl/DsIw
AOh0UPrGHVglxsYXkkajmFuvLCu8bjXodAFOFkOcp4bOnZUl4z+empM09fjJ2gIYYfX0dhYjfUmL
0jWBVxdTbqlp0KQm37PKhm++qp83mH78uPBs6q4o7YzDsEvMxWtekfOza4lMwwSdWwC382hAGffh
vh0xujdUiKm2hlT2fDwjOT0Cl18vqKN8Yt9uhVdy69QY+Jlax4v0jfCHa7lkp8D7NVoT9EYk3b+R
TGSxSQP/jExZdr3QOFsW22n/4LHo0Ai8dyp/5heyD27Vsj4NO2yPS1JOw+7IJkyi/t6Fnd+PF8Nb
Lvx5OFY5bps0tiUNB2kV14hxTSUGIuD7fx0EyySY6qZqT2EGe8SrchM4pTZMBZB15t+4yY0vTzro
u8KgNQZUH+2EYuMeHFILBZtrYF3W3346eS2fcmnQcUwqyv2yN8/fKnllE6Gyn+/ICYvaE2EOKllK
0BjnayfOzNDHnKShf+G9sXNlykI4RMB9/jDVicIKJF2Jd/cnhhabFiDNTtlJSg8xBdQ3a/FsjN3T
Gx7n8D3L8Na8MjGbQ0rdN1nxUqzAHlHKJYFlE697/oxOyOAUxRVc3WuuCmdx65PyvP+BO/Tw8aq9
6zgo2KbLyOQDvMVqI87WnLPwRxd57UidKhm65LUK77gT/W6Mq1MR1pj0obIs/GD+GP00rhdUt66z
XQl3te5G86jNKytA7pCIFhKROyFJeLKKOAZgvUUsx19vZHhYwUgcAXcKojNoVgzD8pbJXNCrrA2C
MtxxgikuSuPt73dF2dh6NLf9P1BbNJslyRtkaAJben+ZOuP5n80ZMgT6fxexTuOMSGKTh3a35BnC
X/LO5I5VfxcyixpDU+G82X1b5m/YulQXMTFjU88L+FaP1IZq8itobp/YdtscxDSm0najcPJsxZDr
D7D+eQsta7kBDDsp14viupk45XBrzPAfHyGExEdFJuwyuwmgYY9WjWXlZc9vNOZ7NAOzGDMoysLY
u1eDBURtBB5U73vU9J8UkzcRE3R1plD8UpLRchXcNFO2D5Q2HhYdBzh650kxsZFMhDn/4WUpjNGx
wWPyut0+XdBBuxV/ezDyg6Jzd3kVYpZuaqx53yFPytnqgPQhn7SSEE+i5BFdlyJAFMURXur5crmw
UTjiaB9/brAuRyf3JcPw87z5+sPE++arG7Qtw6KM9/7Dw5DEc+jYtOpg6SL3V7JCIs/hWGu//R0s
LRNPzujRZJxFfglgpI1xf9suqUpiMyyULUZt0YH96po1IKYq300txxQpQFtFNkD5h2SRw7cZitTu
o+GEbdZTQXKD0Bc/RtMim5gNvxoFk2figmS7fkbvtFb2Ud4UU9K4S6bAk5D8ohMFRHO3YtKZRM+p
Ho/BjpONv8MnriWcV7xkLVInXB9QbBcS+NbmgaisMrks4/06FFI68x7dVSqpieWludoKgDIbWJrD
bSsVUM1yYbWKmCcBCLvW7V8SLw3sUL2k3L01ZlxcXlgfzRJ8WIbO9Vo6UZ6eSnfBwaqkgtekPksK
NTV59hA+vV3LYWGI/r1wuwweoMsp7hNprRwPh2SOOu9Qp3E1PgYTx9UOycxnuHio6Y6k05TUblV6
vvOaDUfQZHamBri/NwVDusxIwbc0JpJTfH3w30hbYhT9NN9tR7mHsFvct7GY+XtKb+z3WLQFmkES
+Jx0/dH3v2EeqfbVtUW7MsDlgMepFJjnLOQ7e0WkB4hmJMIcDvReWp9uHM909e/wTrOYUfM2RD7j
Aaaz0XI+rKYBz/lhlEBEDGApHLbE9tcs4RFnDXKOUm6EpZ0BZsxHouaOml06NMivFnEoRv0B7ZKx
lDoh3lNbMrTu1Q8r9elEXgxKmggkk8ueBI3EZTvr7Bo8hJXlaKkJFF2BtoHuoke8ilWfN++Eil76
IPSZPmnGCpOsWM3aXrXdpX8QplX5yB4qREh9ZzxrBT9kyNLPO/NsJVcVcgIcCoMcFHtSn4uscjzy
UJhOBih6IcwhtOwIUGX9x1opfgyeIemI5KbGaNRW0leRFBa7WE1b4fEldnjm1HwerYn2wx7EitTG
ZpIF8iMTZ+tU9AVBie7VXMXddJjlS9C0XHyMro8F342QHzfO2cqSp+k0vxyVlj6R3erGY+kPJuZB
A5kFg98pFWDVuHJTDVrwuzqTNkBHGZc96ofs1ayiVP1MVLJ+NhJqM6U4ObUcfmT6HT/L+7DyQpgJ
M+qj9HD/R73CTl3lQqsVWp7cDH1R3AwxpUtY7At/EEkL2Jbr7x0CzjWL02BUkqscsiB8MbHQ/TZC
E1+3pPaq5JkmDR8m9JYGbRcfmjqrCQiVduAISL27vVJGCSswQ+oGLB5Bn/43312XDnc8Ig129KLu
CHoZ95VdvQqq4ewdw1AgoL7v+VHqN/xTyLYJGiaCAmfCWQZqoT7qDAV7GK1GWUW6knam1UxGO4SX
DUPZTZkEUrg9/UZXiK+Q8fuHoDB+M6cTZY/D44mw5RADWjre9vQQx/63XlxfC+uySbqe9tNwIRp2
wny0l36SLF88Wn1FMurheiBuz3GvwLhr451CzY8z8hgWNgXSDg7P4QZXmHM9T3vLZOLMC5HmpRqg
dv904Ex+pisjfLk0mxGYv1dFX7zblY2RMsYBsmKH3KCbPrl41zoj0tO8fjJTFb6Fiuuafy/ChKuY
cynnEejKcBlyr29ZK7bKc5QDZhrGVpFYxUisPi+o9+kTMc/4ls623U0zRxrL5NbCEfsVOg/26U1R
tVpMEZxcnaIxPGNrbGBdaomjZ6J4jS538KrTAEgUl5+IKO5llxvVMrfOksi5JWEkYa97dopEkyyW
91/YG8iyNnZ/fHBJySIKlhR8wouc2Ivf35SnOt2FjaO7HEmQ54aICEprPb672PgAaWdwvwl3KFFb
hidgBUV3cH6Hq44wALqHkAb1R+6TfYDlOP400X44a68JiMFT1KMxX7Y4aQzN+Qc0fDVy5p5fgNfX
2AFnVi9m4lNPAP4GKJkrd8F/Yds1HlWGFg4zLu+4v/t4crnq0V7JfDY2OIXITfkxmukftSTxB+Jh
gw1RP+Le0cuS0cYrJvuvbpaqoCoBPrrUPCjCTyke1KjMo7Xsvr2s3Hat1KKmstRfv62sWCOXk5MJ
xkvb6L3Jt7TVyivTOJfeGxNyM4DoCt00RB7hgS+riCnE+Y3gxilla5E8T+I/gRWy1jb14SSSZUl1
3rISpzBHdAsPRG3GiLtF5L5W9hUmfUdfDR1he5Yn3lfsaz4887ODDGI0aKHl3/j4S/YwC/ee1teE
UNYmzXM8ntWAFuitPavmxSNxKI8k34OY0BvmO0zvk7+XKNYdI8mcT8yLgNhZcWS/Wxe7eBrFGi98
f7QNue7bK+G9i3xiR3+VFkva9toTzhYvP6wqqdqSKD24V6AywQxHidFK4QxaF1oNMQKXgfTbloCz
ogenkfoJVjD51/2N9wNiuuMYs5UwSc4g60TVWUb2Lzcb4f2+YC5v99nqzbrdeyx40KkstgnUPjrK
hCE+Pr+gNCv9vFu1bMTu9HfTHezVFGDUIQzJfyIfc541O7KDPOg7XAwwCfX2rYmr9wQU3YaTVRMp
dBEBkUFpAIwIBWuRpMKXHUzO1gKgShEMMEnGqbDnogUmNavtmNLnq8uUxUheDLAlulaFdNW3jxFe
jgyoJRJXusaECn9r79XbyhSq+aQL0A6Ab9yHI16SLi9ElltBJNg3jWULw07TBIoZBZ3uVmpo2Jmz
R55mS6Im7MMOS7ZcQRjAyypuHEeJ4TqHs/+IWzqECVlVOR4XUIhlcdZRw+yKaVsbpZdQct+AiuR0
4lU9PAoiaAJyCONz4sJxJYgaL/cJXjeRFsV7bD7jYUaoOYxIwCVb4ARGixqLaIqm95Djmg49OnwO
s9jT8ghd7wACtjQeti07505MddNGn4/lxoI5FjvUmSYTUTDbL2hC0ta6qXMQfL+VXADJ1Fc56yNR
ptxoMZssxtS/g0AZLsJAyV9ebt/hRxN+hYagf6LnSN/vpBGl5qMonXgeadlhAJDfk8T7Js5qAqTK
jHNz/ayPR23ApiJ9/6TdvaJV8AzEoYmOM8lF6Vr9UQ9ZYx8nrD8RNcmOKtwJCjd/0fGobwg3QagR
0bNGRJ5nZmA25tqf3ThV07nc7DnFnkYNGTTxwwurj91eTzWIE8Fg+eMqvlp8IyucHFnLSEqW4yPz
uDlhrlktac46kZPLqfD+n3H/DYKub4VVkV1JRrKkru3eroMKQfOTySSS+lTQoXQRT0pmKcpqUo3V
3JG5sh1HZoWbd0N+b04UMjjlaOK8oXfYgyGo6CXl1R2kmT7WAXfdTmrBGcAJ3KivgYrPLjdbkkge
Y86Q+LxptZfXyuxjdJNv36d785SrNARTktTbPD5op66JDmHaoaJ+dqeEDjKkZZJ0ZKOe8CuEXkIU
UroXvFgD4itZHhNLdtnCVHKsx78NjhFWx+oJID9QhLtLGH/n+1FcU2FNcxmDsHgnjGyHGgy+KjqR
NWob4Ij7OuVE92UDbtOaxD/AFvu8bGoWnNqPjKrOtc27thIL+mrOZ6JV3GJ1h6A7oG5nm+kLZSEo
mhSo+Cnkyil6cRt+P2LM1QKPFBeZedVCIWcv9oFyv5GX4PTmQPqX3S6iMDOg4LAsZU1qquYGyfCW
n1EBy2VDfGfRw/GOFgd7RFPpreF7MqpGvV92UeMNy8+EFfGA2j8aXa8VrASUT5V28VAkoGIqt2PL
UEYeKxLZyOMv2v8Tw1eZqDpJRTG91FdncqL+9B9ccAWbP3+AYVkZ8TUw5JB3f7Qa8bKvQHePAeAJ
ImgSXiPr38+tAp0GOKwOyjgjjAJT1n/tL9F77MOHqqX6R9Yxe0UDq3RVg8JcP94FtTZ+0A8yWyNE
CEsL1Cq0Jt0AR5dzmgjNSiogYXt50iI1n5rszybpgSuGmA35QqEt35/eHcc9KKftQCec97s2h+pC
C419ENssIHhrI56Uk0dsdBfd6UCUYTxX/oL8SI9BSadO/hhUWfefT1V/36DN8qpfgIiGTikGGQjv
uMlpfNZzMzHPdpUSWxIpO63ToJrhuke+wus43bWqgZJzzerUPzreLORBfacdAHjPW3+XnXlebabp
l4Y1vaM04a5WpRWQXvcWH9Qc3x4H7dU8w3rR8JTp3N3KSYZheVEgORmN1L7e1Ra9g7XQ/8DPZqEy
o/1MN7Mui2mSZlpwHfe9p6LWoU3F+DP19VSI1+3K/ieNNU6hywzJnBRK0AFucZD0SE46osAq6pG7
ZY6FK8PtH58/7w9CkuxSeHBW/BckiobX+ugib6fvE4dQOi3SBtkrvfLOyPbtlHk1wNvrE6xTqP9C
yG5nirsqIoCBdMWntCf293+YDAY/AdBxEYekMCgYGpV5H8EbsfmLOCym+PUfs2AJVOdQMGTwvzzj
vPbpY5k1Vwdh6tVEU16oQEr/QqTQfFI3zh5ysdxgTQ2rH59rxDV/VxeIUqPtPOyAxyJxpwN/pEYH
raUvTaFlMUplFUG3xpIMfx2zEiAvu/bmOsKW07TTjoF1wH5rBVLVjfUD85Zk8+tcQk1P0T4LYitB
nYIu1JznQo1ct/5I1C7ere4muS+0BLoZPP0FIq7cuciCuuv5iRx6u3gImQhFH9mBhYMz70QZLidX
wTPZM8hlyV88JIXHDSWtlLRHk2WhN3dh+qfsr9zxksb4gudqghZQbQreFvA5iOuslALkQFtu+AQV
t61zKFSgaNMaLfXCyJvni24cuE+pvGHRAemo+/P4x26MPZhJQTBGIvKld2+LarjnNIxR2aES9Yzj
u2NLXais9fhHvfd2bTrqsMa29ogfEvvTliZ2oxxzkbB7axbhOYSOJz+pnPMBDpO1wb+ypBoL6LLU
QKfcdInE184A7vC/bWXarpDvGAJCwF9vs8e1X00HFWf/2OkZsTiYCsKSRsrTNTvIulJ1ZXY+0SRB
+guZ2FRP5vGgtswVYZrwmLiJMee7RUwQhY7tWkPkGDdTsc+p//iGPToS+vauy0fQwfxCgXK3pf+F
rpcpfcNbSJaKqdFx6h0JIG8EeejrGvVsXjVQwu7Iy0h2EO8m4C35BiRtmsJoGTjKVPf/PAr9ns6T
ODiXry8MW4I31EdUOcfzn+tYuNC5TAzAe8oKHnsF9UtDnEogHgb3pETFUou4E5SWFUWP8cNc2Cxw
xsMjlc0cAVIZMqWxCMVczz/TU2okHPbm0JipH3NOQZJV8Bp5AZuOz8fAKfg34yd+NbrpEitc2BmQ
Fe6KGVu6nBVxCQfmOhIiwBNWffSj1VQy/xXOhjXgjfCPdmD3uu6uQUJXCBLDoSK8leTfCxvrqTqT
Zp7vfhuXRXXFCdZ8JnnKo1843E5roXpe5EBssZi2WJ0fEjkOdrrkmcSq2K/H3ltV4uwcMd9dGjqY
A9FrNFZPk5/nYUNjRem/zgyd67vIZO7DNw7RPLhjXqgIKxKB2w90K4sCfYEHD8VzQ3+ExJDGf2Pe
fBO9LoeY+H7UxeobKvgns1wsWrRToY/MpyVJ4HGGc95T4bvjBiD+LVfUGZ0m3RNYdE8ze0humFQ6
hpDdMRoexD9Gi6K4lp+gRvK57tSlH8zqvaF4FX/Cm2GDn66jkjc6fZBambD/m9/mhxIWWW4d8mC6
17JJWwOSNSsEq1kY4jeS0oUlX3fs72o3krFHmRL8iXJSc3jCTATLRBw8i6P0HRf0xvahkCEpsIYT
VMj/KqFFbFBpUYdnZObuXZNj+Dwoe4FNdlzk7fm8hEQ5L6W/9SbBjxUOe6gdbKmwsAdBOfpPn/k8
GcXHZQ1ysX/n3QJzXPgg/YMqwxVM4hAIeOKe8fhEXV9hR59vMy06w9h9ZP/RCfOFASw80dhpqijI
a/5p+8zRMs5p5/MTWQD9AoNDNF3qKPflZc1vGwa7fThkK26YD7mUypaBNyvLjzz394pc+LkOIpcO
67X7nRB+gyBsiwQ+d9RCG/nQPKNVUWO9s2aZV6cJS1Z8TbFM9I03+1ByH4GKD2FFkMY/N7Tjaw9e
WpkbHwfAxc+TJscGG9nfxMeWDhs/OPJRr6uAKlodXz83rOsOcQ595XXdmvxBSzkqXbM86tklk2wu
0VPenK7XRRjb/fz29qtdj7JfGyI/taxPxLpiWWisybMw4oUipiBx3mhrye5auxWY+stswMLSpr1j
dy5CuP8IvF+e/7Vlb3hcNPG6HrIQ36qvbUNyuc9/gtjlhgGHvGc90xPA4Y0rOsQ2SzcT8F8b80RB
5O0ggsgHtU5ZTC24kIYAXONhrBEdFnAVBrlQxI0lwUl4j/mYiAw6SISpiU+efZkefv+DmkP4CvB/
542HgWje7Y3hg04eph48VnV2ZG+JfWt7nObG4U8Q3eCNMvWsY2Ojqwv/wF8kytHiHxo+LnHqDSrB
ebBCOpqBmS0SiHfWkvjGhSZHMUSne1D1t4oO5rU7fPsM031obNEM9/0rhjBqKpK4x/XA8kk2kgyC
B64MFa7n4gtmznRmYnYMczbYbDUSRAhfVw10zPee+MIYmj3WR8qR2HoJdK1PqNSKsIT1SYrsz3+c
7H+y1d9jGExCB6MlUkLuRcvupBO4/7i2PRzFfsP8bRXnMzi9DJ8PXdQpEPfzPcUWbWKga/BrR4zA
AltESccPkfv4xDPrNrRU8PeWYaH4lRAkNpB2HUIVVHapQJ7/QET83US908OqZN7/qKQnVHZ97Qsc
GvEF2CvHDs1+2GBGyGjAMiobHxUccSIld1ir2e0w9EEkPk/aIk19KAEDor3wVK/HfgCzP9sFYueq
Q7ULBztHMM3KQ2WgD8N/jMWoXID4amARL3tfVOADf2Ri5PZVW/OaKIBDFqVdrqNgHivf7Kflcywd
0q8l6tP49ZVTtL+GQyj/8pFqHru03PY6JcrIT8FMtYRrYVqaMj/GyHtsGBPrAZZzpiBy0bhxNYDz
NEr/CsdTb7pO2yHqjp57NeJsKWd+ZzUbtTcE5AixrPvH9MvVpqlcDAztE6BbnWD1vQ7+0qsmbvWk
Tq9YcstXXEY3PaDieU+LOfbRDzEu9PAgrYYoBObJVz4cwZqZatY+D9fzRu2jkpBdtm3NsTTX24HK
F41YlKl/LLbbHVP3PsDpUKnvd/7zgx+9BctB0TuYP9jnyAM7p2v6aDxTJttjdm9V4kdDdDitjzJo
9r2fV08ZvHhKMbu0T9oWE2IFUMbeYXNsqpuCjlkYbyIe6pDhnWlQbMZGFGBYNzHGwVLIpsOsci6E
vMV75dr0JVgGT3doKd9sLXCSA4J5lM7TVA7+fMGUnRWXorJ5RdV4t/dgZeHF0YNKymLj1cE4IkVU
ONeH2PIPkhK4OtJK4O0i2MuofCdSiGs7C8nY5Rb8vmTxXADp3vAVNLLBjRqSLqRxFgzeIWk1bp7l
Vd7qlZBfeOiwAJ8Kw1FjeeQ7VXJKhyINVWfNXrW63MUJbiabyv50w3MHG7loLjJRfmEhLeor5/L/
UKOOdEOVoTKIc8z54h7eug+1sgCVKmULPEhe6rAk25e/cxaAbvEME2XC96geP7mN/GW0XsGIyEJS
kF+9zawq/RMo7ECr1dxi6ZBSYnHQiptrGygW02kpUlmO5sq5KVnmrmNekIKYx0BVvSnOZrKClAWM
s2z196rrpmdzsGEMPp8oe13oMNrn0hsMiKln6MttdzyHVCBT6ldbV26L8uni/LSxcSBSj742C6K4
dVB7gMawxY2jqmovI49rQ8nA02j/aDEd95t8p3DMLx3SCyVtgqUsq4DVEL5jbggFSXAP5DTjp2+I
OIEluRfoITNJHrZg8Pdc1kPLhHS8MqOoM81zRhlvoikiKKMP8fzFeniXIMwZ4ppm4wDFVzNvd+U2
QSb4r8qb8/wk9mDwgIebLmsuSqMmdM98iCdjsQU6Dsef5f1fYXhz1ipY8BSgIQZUbB+Yognmb3H8
5B/l8lsGWCu4RHZ9GQ4TvPrXjSo6WEnl7lhfSn+EV5LkiQbx4G3MBSGitZWVniuc5nsOgwIKLRiL
cdxDF92kXZE1ae3YxhnnvWvo/nNHlSo37E5ILS5jEedtO4XiWeK2HM4Qcy2jiQ4PDUs54FZ8lFg9
qc+FKQw3T4aH4O0nFNneBkjTpjPhuGTfjAZZcvVFm6Y0yXx92vzdMUtScJ4Qo0T2JojOVuDUhrYe
CKWfJbevNKPTA2J5TgftyjDUXU/+1D8FrNQP0Wrbn7OZLyUzN5esOcjo84tR6mLbmc2CNPjr2mRd
a7OKL6giX52sc5rMnlrrmynHCunBRGniM1t5oWrSZIFUOlBPenU/Pa2fvchpbCjJlmULR/A5lQ9A
BUEOaEXeLTjqS+m8i1QfPThxoSCaOHb1nsIzQXLAn2WFs0Us+Pny94+NKX+jPCX3ax45i+/aBWKT
sEhZNknSmaqpHUlhfZB3ba12CBTgYG6O1REduIZvWoVJKVE5nNMBpGbwE8qoRo1IdEVs9vanf6fI
1E8PvMbGrwazi1hQ7Kg6ud/Veoa78hsY3GLQbdVGVQ7K+J94OPdctPhD9gsGGv3ReED3DTctc4BO
Vw49X0GKrYhsH1LN/TFHCxRyjCfKFh4lu5VMrvKnelaW+OVDCFfY5oT7hPfkfvsjf1Ri2s2T6r9C
p3qrN0fOEfBlqP9snHqkBlO6OlipJLHgdTsew9Eu5IERiwpP9wIuN3a9Aecu1u0Vd281w/xOPxKv
oeXyEG2Y+JSDxm+iBRVPJAlUCjRYaRwcilJYCdps/lSypdMvtjkf8yyTqP5GeLzpHwpRvY3T9OC0
pV95mutLkVWmREBOiHD8PN1Lz+cG1MI6gBNGWe4801l2pyTIhDpxyRAbPsd3LBieW9l3csYQjY3O
0DRNxWxLtSxPrnWDkDfOK3o55oDgoc7o1RQEgldCmWcQR0ElPEeZ1JX2dHDT/7w3l5ZEhEbSqggF
XTLDeMttQtJ4DsPL+fyYGNbfVEIoMzFt9LyaZ+joaiAwMJXfYl0R2wXBdRibqKR5MNsLVSSpNKmE
XuZZQS9P/eWZ7KRqeoIQ8kugytU2vi9QyCQNvL2OosU2EP7s0qT1MmYNljZ5M1bVuGtr1m56Lfjz
Q4vDRCR8JVU12n7lkrwjuR/k4ksgiBxLSa6JDUx8jn03jUyIM/uZswGGsdfKyiySWcZLdpFmzmv9
MlutaaqixMxx2wTbijaSBVDC+EWeUS4ZwhAKSYFFAnU/qkMiCwzUAmIwQQiN58cniCJNGjiap9ZP
65d2dm/0ygzn+4UWwYbrNFcfH3XyS/I8+JBsgIdBS/Mc0d/eiZZ3Mj3FBUl5GCBHh2bU9T0eRzWo
3LTfPIKnvHhIUvxZcr8ZwVC6O7z/Vy8j0y15Hj91nVUAwrm5JhYEI9U1UCdZTYwES74TNhrGe7pk
G7WUa6WQaY1z2Svev4irf6dtzuLUj4Uo7YUMZyH2k6r894GswJojRqccnuHVq6Xr5Fos+GWpYwfV
yRbVU8RWKHzWVUp3L00wEus8L0y7ghANG6rbQL6eAu6T1/zZduU6BffPh/xboQcxFZsx4iWbhv4C
as7RdkEPdV4TysJYmR3R5j8/fGG5xeunlZZvwaib5DBTbhHxDe3fREe/+NRj6g+ejHoGh3ucYY1C
CJIMOEbWLq8Xx/s0MJOZnHISoevbhtwWmBjOCprJl0YJ4iDPrIbHYvGYgOCUN/r43r7KUPCDVu+1
oo5cjUFoDow5W/8xQSLgk5rpgZJfFnAsTwCgSC59OwxQRXMN4/BkUagDkgXvbdZ6zuX9F57AYJhP
Z1qRdA6aXVt3ZslqQ3UZCMV+js0cifZeSx6fiHJIQ+HmnBO7xE2t8nld6Bu1qD/5Hwbkcz9+WUYx
J2rkKce6bVPhz5imD8Ri4lkJMrrr7nru8YYIOQ39p+4Ur2f78WwUPhexPT3xZjVjPbQycAg8Ahcb
1boFKAYnUYJmzAQy3ki9e8Zqn7mzdOo63ZX1xL4dXxqQrFzQObq9X1QHgMqySZQpPCYtQhXrA/RT
6TvgXK7dnnywEBBGeA2soQ9iLD6Wd6dskj5MJPLASQy9TZof1keozcnoZPOEhZKbvk8n62wLOE3P
SAawOu5z7xcKheA8xhbr60ZVKs6TVN2oXiWt4+rWF4AtCEGY42Su2PcQv7uqKNjueEoPA6I6eRR2
bysR2qi9kLWrBljySbJTrOzj7JkQIdC7AELK2kIOhGUHtPr7CeomG32pg4eMkIJsLiyVz1Mybzxz
KQQR1kVlkMB4gmU0wCfaE2zmKkAQGkWxdt9nzugdhWHk6XpPdIaCiuCj6bz4bOAYsKOYcAE4uB6X
pfVix7jj4c3TufRpFgakljfvMXKvXxpjoRbuvUl+ABlpHpHSsso8y+fnsKq2QTAM+842h5KwZG39
TaO2jdPbtUVxLHm3lqxO/ICrEm1qjv/3CQ1sxlqyuJsU1VUbzk4FKUx6Ca1D0DffiDg9MhhF7hkE
XzzgC+YRhsj5WdElH7b/1DpjIBLL4txbkK2lEc93q/LoNiqpfXxQfCpNCfudyw2eMg3Xw++CjoCT
lQJNFnTeJLWSoNErR/4p6oxTH624MFTNKxWyMhbsJ8ofL0lzKwi0Bt2FqrCFrgsg0Yk92lwbxUUA
H2nGOG//4C6CnUzeavC4kh6dPrYKepPbBw5y9LCv+njFnXInias1BVzYdSOnlhIRRxDRLWyk3lkm
z1ceH+wuXUjkhmffk+/mSoR8+8dR8Z//c7ItYMS1SVLT6O927N4QPO4DnK4xfj8gy6uI26XvBaNO
tJzBEAxSnmh35qQ7ug5jc8aYUW+J6CZs+aRAlyheGNTMEZcwTSxyFKoal9SOWMUtRjRcUaMs9LKP
KNsiWzhxxWfut1tP+lg9uRz8ogNHVylARsC4IiwvF5qjeY3uRrIp6Ibh0JcBFdq2RFCxt/EZbM69
3y70gxWAETdQ9qydHdP/36KGLz99wei+tERLblJUFpl+u9PfGPenPg6F6PAhGrfxtjb2ujbuaSyM
+icJZs3t1Jyqopw7ECQhuZYEKx0H9QQC7pTiWi63Qu/1v+U/Lpvv091IjZF2McCAKIaSeFUwBjyu
deDVSljsGYzL6IjsxDZdXMkpcJDwKa1hAd4k+K4B5nBfSH6CXxVBxLJ5saspC9su5ltNMpi5m9la
W+gW8L+d5jQIb81FKduPROXDXIw7OqlvIsLNWqLsW2mkHI2HyBVBK354RTx+drohADefY+pWUIrV
CujDGt6a778Y0R76up82G+tQokYUrImEm4TYyzzMF1N/EKNF0RiOiV1YYgIqbbw8VtW3+a9PVucl
xiKWEcDL1zbaV6fmsnUJ4XLbkgkSqgN4zoHS/+ZUrero9GnywcC9ZgSZTKltwCAGefJnXYKePede
ja04ycLrKwVMxZCxZDqmktaHXv6rLSpR3KcwrdinOLYZ22ukxkWURJaxaNP6tHKuIjRFd1RCZfH3
WFxpnnXjSLjhJffTgMHsIvDdEjiisP9tF6zDY9SUL/NG5Nf1f0xJRwxBWBTgunUstDJUkrE70sZF
25EzeNtbcIZM+ARmP75S13cz6ME9Cf5dpHQjkWe4u/7fUNWelRCyPQANlNprY6oRAfI2jAo+BMSz
Lhkx+JGVfPLOOKkuJjgdUHp0aTlhJ6uuibQ2muU9UPATEeKUPxqBVDib4T2lMi3ihYZGboc3AY2m
O5B7LfgtBavPt3MmThkhVKogpZZYnTxlmbUIrwXjBSApStfZgy5Ps9aI9Hftuoj3zshcXFYZ2C4O
Rs//NBhiRAXIkz0qRsYlNvLx9henmOeQj3Z2cnnxcAk0W698qCf3F6MoYUKMMwLkuqUUO4bz78PJ
y7AIhlEXHgvHCQLJTJCKMbKpZuJk43zxxOVxUxPJdvpxrHtPBw+9UAd165hLX5mY/QS/FWec82V4
i+vn70c002A2a44t9xwwIqm+/e/4cDDSBeCjZOvmhig0hOErsXrVfK1TdpZNDon+J6epn9mkf+sY
wyz0W3b9crigzg+ko9AW2AZAegvMa3aoMwTIlaNa6EuWuAzQGe2M5Nem6BNn5NSCulYX888P8waW
P6LFmejcR90jYbTlTYKkc0OIjlsULg+tB18nZSqqKQem/aU+fX2VAmPhk3OaAcJu+uUBt0JyieOT
q/R0B8lZ8PfBE3BA9Fyf6k0j2ds2oxpE2Wpg8nJd/tDFCDIr+qyztgo0jW1oYxP+kU/fUUUn5U18
nmr3mrPvglaVei7LbtFRfmz9dSutiF23/KJ2Kht10ELrWBZ4NIkybYF7a2z+WNt1xbU02QjFOzfT
wWJkRe8vJkgRZUlhBbS3JoJQNmDfNil/HjvELuPuyyJ/Lf4x5t7+/3sNgMJNLMqCfjUOXuc+3yz/
LQeJVKVF2xiTQscaOgNwFhlC9mBdsN6b38vl06dDjkOIVGW5EBC67JNgWLV8DWU8tkOS2zGRJkbu
2Gyymjl7M3zrRsRtMLKyExDb3wzuKx3pfuBEFhD6IYZVfulikjLWg5tRXRHqKt2yUZ751iEPoTQv
tB9K9Gy8hRvLijXihCZpVHBQXx1guhh4nKxol3jTSSfm8a74gS5qO5J6SyQOdIgI0Wjd8iVyCha4
pHC0p0k+0iAJAIDSIOPVBxPoOMbNeqmnEn6y5y4RszKYA9ga2W8fBxacchYHIK7UUm3taSyoGTsP
JjaVPwsqgf7EqM8HS8YrnoznGcob1eMas6FKTC8cZBkdoVhuD2BFDNYWCOrDJf/fOFaOFpx11mQc
4F+1opoQq9d3F4VJliF3VVx7QwUl9ItGNqlaISmSCRig+XFUMjGQow5MxKN7EbvGhDxUzKPLuqMT
dHMk8eWwJj6kJFyi7YvuJPbbuuWwuZbKaS/4nJzBJCWNyRQ/sBrlKysbZQ+RwxrLol22HxcQqgTx
ZKPvtol1t9VYnkKY1uAc+pO8h3l+x6r2EbGyvg5tcFGtEKntM9nlxEcYf9qQ0HWvtSdWLGpRE0wa
OadypgKjuaWDpvr8lRVNvIAyPjoaDPGBHxlatpZ+z0vZABmsXgF8scU0FLh/eLQX3IWPYQsMiFkG
0o+8dNaseEwcNRSfpwl+rcVFkTVYCm/LzXsRPHYYFIIR4k6i5pdKVsEB3wu1pDvTRBUejCEE2GzH
OrM0Dzbgl5cj1+XOyRyENKRzLfPYf21pM+BCh4fsKvj2cvD5MGRVAmUZV8oEeOAmXkieFNnhQ28X
pkjTGKg/gMy66vjoLF6NQ40imNrkbSg7aXbU07um0q0VtZBlP/1WFs8Z12S9VbOnxRXK7AAN4SH6
CZqxZ2pdq/2zzdAQkafe2ImXlu3YnfcsZHEPhlMMiD7NwT6ZKxpNEI29AazikLSQSKFFAErsI3P1
eRgXpSnDIfBvRhepLaohay18bGgEKAfgOJ3+S+Stll841RxLSIrb/aJliHfFTjcIr1mU3px8dUuv
61/YbNDZcxrXRS4h3FZkFjGW5f98vvT3nulZhNg5hMV/b3F4LA2wTf8Zh3/Vrvv9CF6Ja3NZDqI1
E97tLfSserw9P/K/y11uMaJozz7PhM1aWyoyBxE/bjuqqcc2OZJrIwbrJVyw98Zl37VQxNDJBDYf
68TZVR55+vihjhe/zU8Jh7C1LcR0QyQ3x7lMD9t4gEHdI/fn4P7a/2HbODY9cHP6/lGgBWUqfn/2
z4H7SB4HnCZExccTuPWoupDsxdGgYPEvP2IYy23kyX2mD/GUWOyFQzooALos4jdFprJ1S5qmBT7X
qMAx9RIk49eFyhYN26GnBWCyKm28A2X2b/kV5odTgUzk9ikVo7FzvvxRalqmNTTG1mD1Tc+TlV4Q
KgAUGPOFx38yalsRPhSpGizqB2PpG7OKTt6V/0Al8UV84spe/3JhdbtyI8jvnWUW3Yve1dLbzR2e
yOOJDp2dJeRQSqJzyEVyT+IlA8+UE0j2TCQ/0GyImhqGoX6ltrhx3PwQ9EEwsMZXYN/BeyaVkZG3
6mxE1jXbwtcnv1MXJLnzbnBZVA/I3yCouSEWVTDCAvFkipoaOfpDRZxzYcRHP4OEYOWyPK6pgxmK
RgXuvxR8e9YIPaC4+zubmY6LUCHB2hIkQXkuGhODTCsjGt51u6qxrm7iyomGgg1d1KR2xiKPR8Wq
VPlsSo62748X5H8sT17iyvVPaTP7KFX5Oibm+TI0gZUFa6TEa5eXBKZiegVjm/8IFA/Vtkrhzrcj
DcZXGP0rqM0+qBclm3+gDGfQNe1Nu/pjHapTWsHvIV2+da30lLi7XWNYHu2X1MdgM/j46PSzfBbG
yFWfnjgk2at5yIF5gIgDCGJeDdL6Qgzm2LgsxGWEsmzlZaVOPSFsKC0K7q87J/4t/vGBP6YVVtag
5hpN0CYv8X5xBpXXYw9PpKTVLbufgdm8VUUajEDvGHXign8gemxKA02BBOSuUw1Ob6KspsXj8mDK
6Z44HnA1TQApUKOAR5gf5cjU/6jfHJpAFEHbo8R+wHV8SvwSfx623ul4OrVJx9NidUqQeu+8LvzY
O0JRCjc2njWUs1FqQgtznKWxeN59mSjjlKGmm8P0udA8Vbu/RA+46Z1MLQFC0vUyNz+RYG0rhQXe
ouI1eziTdihDR9uf19roizC67FxlMldekoTJGD2fJZfdJXar/1fh5Ys8ZdUn1iYeahjaOuTs95gk
NLRmg7ubRQUwBi3odLOCzCJRMwRTFm7MN1+Z0biTl7g+goWuqaU7wGy1l21V4KCIxcTXyK6jia/S
Zf1xdhBcw0+f25o71nZx0XYgoebYEQ+X2sUO09d9D2pQYdOrtDbu/wbiWQZ+VnTp2b4dABrNMYfW
POromUnpniLWuo7ZCrjFpfn0i/JEm3n+kHOSnLEyhUCmRwB8wp/8upYVYv1lPDspALo8majDq31A
r2H7AiAt/wAKQaPZiW19i/RMhU+WDGRPNZ2Llcaldbod176A4gDY87JiupoduOFOYQcr7Jv683dn
iFy3t0g9mLDf6T6ib1FUDT1GA9B18SA8VNYXPVpZUijs52lE9A3uWMAp6nzjNLPRBGSZ8MvJss7k
FxkG9YBWH9xipxV0jl4dimJGoVhbavabMxQnzCKzncLCk3d1fWS0qYBi7SvHbsgI9atTzhPaL1Rl
4FCxdhUYk/CkA2smdodu0Y6IAtPcMzjrRuSUdRRnF5d+NqST2IFXZ2D6LYuvchCx+zJ0IkojZopu
qSQcnWs349lRP8U0QfYJ/TEYNBidCjMaNnoFZQM6EkUR3UFV4IOY74X0DkeGPqrpvcEs+1SgkhrD
Eski6wuzfBxyNNRqXCQHw3P+w8oMbf+BvyYnRrDUpALUWP9eFXtPL52mznskBx9c+X/QmovNJMv5
FcJELLmwVieTSVHS9BPG0MDyCwqXRhP2mm5qBUgggg/qCnGY2yUcGjMP2STdX13U3qfA10c2wXql
94zV/tw6YyfhP/Iv34hvS2imWq15qvw1Ps+c0IhiLP0rqGWyJjRZyGO2iD7t69bkwEH1h62dTdte
uX2gfpdOHJGeWL6pKVZZ1ZkSX2XxTiBsA5xWtNCG6gocxQ/n+jtDWoTXB2M6yMvrSIxUd9wxV9Ho
YcCTPKUJTpiVIGAHKgnaCyXGGvdj4ObEsoLWhRG4JvCrUkCkAGn40+P77le5QsRc5ozlea3i9J2+
G8FVdNTAEP+FFugWZlxx5SLlqQO1Jz4lQcx8s9ZxYVHyHGM3aZ88TJ9/JjFi/cB+RGLwL26IENdL
swHEdGqYs0QSR2g8RMPzkRelgxzifoAcwkBOEOiqxJGOc2t6hMXPbMDBhz024MlTFfGV9iOQm2VU
dIUbp8YbqTFMyHzKigvGxTJUbtYfQGUIdAtPvr771S9ioLk3z/Kvt+/PBbzalWGeiq7KRokriFWx
7bZ6PFYf7PoSR+BoJ+03ZI3zZaOmpL3kNJdI9ZVTSVotJPWHtbpz2mF0jZkOaqdXXxZlEfs73rFN
ma7KSzFs2pDitfyikY2/+iNppZozhHqjzE5G3/Ab/wh7P/DP/z2ADGpIiLPuOfWz4asv13J5vjNq
e4Mokq4bW9sN+ivuLEs2tGzxTux/5jgo6lxmz6eDJ0Cw/CICSI5cnh1XjlixEkwM0k8CPdEG5VMO
gLH+5Z5787cDuLGzphkKyMg7JeBg8sRyq1ZVcfuxFViIRRdyVNe1stvkLn/zfE8o6DEBJPS64VWN
lY9IkcB358W+Z5tKNLBVnAKocStgvLUeEgRJ2zPxK9VoKvmI57IXOKjTzWLIfulxF1GqQika6nG1
BcFVs1jaU04ChQtKigZ5S5gjpsOnee+KhRy843YqBOsmsIWyTnYj6fnPFsEwMIx184uKcCxaAQQj
1+65wgt9VrjVP59whaWUej01BmJYM5SF4cked6FikwXKuNAtsILwbaBQZzWHCFAmmqW2bIeNyO6w
wqLQa8jNGVsdHLfpwvBRKmyLemoKSwZH6jZLASnlnJIwefSlkc91fvgb9nHFAkLhowyFJZCya11T
b8PcvncwmbjGHyqsuGMn09qCh8HAa5GK6EaDA9T5uz9E5wvRdRT1iTMLf2SKODf4XET3U4gaWXRK
nqlY/KPpOoaTI4xLB/FqrSS42W1WhzA9jnvUIzfgNMti2nptraAaelzYXkVs3k3X6zveGVFumW5E
yT1PS/e9d8pR13iAhxQBr/7driGkQRe1pq0gpj1mHfTGzZ8JSd2YEZdYLJ/gQnZbi+mH5F6epkRn
UH4WdvjfNghY8kylX0oued/rbbUa+TYhDrKrBeZJgUo5IgiEIsrCTmc4UQJWBlUK4Q40d2jeJjBw
nzIAEajqdpG3/RJVFkPOVqiuHRnp8JD6ncwMgGXYHvM5g94QJtn/4fb4mQVcD4obmhmmxOlbJLlp
FLgXiENN53A3yURo0c4mgGHBpy1ve7TR3FgUkE/6JMUGImqismiOVzbaPS+SoGY4ee4KgfmM8/+m
vNAowJlt242BalL491OXu3JkL7ta0mHkikvwVGAq65BX93u3BLu8m5SZ0V+Wvek19Di9Bhuz0or6
ohht7SlLVnloFzxI/nes4AtJ9JIMjhS8BaUoGq88a648V4TpXdq+L0RyDuGednYTm3KuauvOWwh7
HAn39IijzICVaCxhXrFS10ok4gDMZN+Zhuun8riff/I6cVXJkLyWP4ycygGwI6m2ldM5c/6bssEL
SAZESDDUeWqJJgdvXkOcXl/CLwPHUrLVqMPVZU+YhbcIKKpLTDvWEwPvHuRAvHu4FQHaU/0Tgm37
S8Z7F4ypPKgNfXutf1t6wpj4z8ppOUBEZq1GW0eyFO6dbUb2W2SLC3T5/CVZLsA/6KSRfeMSnRBI
jgJMvk95Cpwf5F9V3nMyXufS4fqNCHCVqVQilgDE5VsCTHEshKb9bIYXJxm0Lta0DYQH4aA4wiX5
T51Dbm8qopBjCrIiUNGw1lnmXO80PHisZRnuTWXNegWGfMIzJv0v/s2NLyyxSQYWS3Fn++HiEqZe
9YBtm0CEKyPCJgnWJNDfWf4xEAUOFRyOZkd6/WImkPx1uUKD1ZXbww5wZQWpfFXn1eTQA4rjKSrJ
k5ywNsbLSPI7xpHPdU7Zbv5THrt7LaFyW1kFSfEMA1gUTuhJJPirk9fjYp4smEkb93xOnmLHEhgD
H5kZ0mKVJtwM2LrsL+Kb2TS9IvWBT1X6oMc7avEojWCVp/ayXmP8/F8y1+BnxhzUR++oTGvRMPm1
VFxWQ4U5d9IeQMSWcJmXVAwuxQpTRyqkzgjVxpovN/Q59/bdEJESKGel59ZaD/LTzUrrWwcAKuTK
bCNxnvdoHEpExtsUO2DzaWV6hahCpUv3zNTBc2zsSuJNwiKRdMQLcI5HzEBQtEsb/akCFlzhwzl+
8f5zg0e2uaqjpRACDrg9p7RkE09oKtkj3j1NHz7rgJ1jt1oJ0HJVz0oEJcRbxhTVLihK0dJbQcX6
W/HWufCpborjxVu4Tj+FYUP0exJz3t/jg1LHO8R5A1bJoJcExnx4mrr/lbRiMsL4Lb1nF4pnQ6LR
f9CmcebMENGXuNEift9YTfquUy0XAMbkbd4T7B+7+Pe/emg8gzEEEr4JqksjNVll6pEi0MLmvUic
HF5zd0O3lGkOslxtt/FcTG4tMB6En+rqISJ2skZU+GV6CoXuOtmO8rjrO1vs+QXWASwBWX9RQPt2
qb7vXDPNNvaw/gHPh+zGeqIU/t2UHjH/xSAnL2EardfNR/lLOkrMCqKJOVepU4P4VsOb9higCfl4
ZZMCvvF7uUVotlWAq2lT075+saL7nJTeeWzl7oH+YdTMRWPM6tbAMx8y7dATKOC1g0cmohtnejoB
3KkkbHagsjlNYuwgmAuJHnH9cj5dCiOaVlnMU/U3NS9sfoL09LEUObFQFETK6U0PwpUiuSx0l+/w
1Y6/7PpC+pUFwXicoiTW95aqFSnjzK2LqpgR8El6HTxo+kPrg5AEoWFgixkiyOITfASY1B3Z3BhV
cKI0rxn6Pq2157Z/JtHL6ghg/ZPMUv00bGdhnPVoEhXf/7kOorz+ov4fEsDGjyW7+hWaYT3SA6pc
ax5G0h9Zyuc/SL6WKzVFnODe0M64n3q9h4rCHz/Rqxxp+MDdBhM2c2p1hajmGlpl5o7oMW3h6Mro
OhkAyG6gDaH2yM4yobzzUMxOp9JdM1mstQQ3cNyzR/o9/ppM8ze+4j1w38yEA60aVuoeJzLk3Kfv
ajTAzlR5NOvagZZm7aSNOxA+REtNe2a1aV7jl5l2OGpLF2Y/WdvoItGwqizF6Ny8GoP9rUuJPBuk
0X7ZULfARHH7zxwCYiVcT9wkTiUzJ3ONkyXWePE2kQoMyzKFSr97/irAKnJHPd76gCsgwsh68mks
sLtM+wY+wXiOjBpjObJajrKRa6LGSE3ow7r7rYl0uHnYvZb7PVzNzIGcA/UqLjO27kl984CAA22k
QcxQPzC3lEB/JHptuuPTO4cqaT3IUu5gBAkeOK0m1V7hWtHDYoi8QkrBabUJt3Ue7smvLS+hvwrf
XuJmz/iEKa+1S05FyPXYbR6Puh21ItK6ZXfxhNvYkiH6WN6nEkWx65tZ23vNqSYm6505F6gD4m9Q
bdv/mFsrBJt/zkO9BAKbrtNVoij8I4lISH27DDQcWK6eAp7HtDO56FFhCQgz+d3gahoWCuufPRe7
3oWyp1yuh2Ab7Zhmisj1VX1MYBKcAdxgrMEnpZAcgbz/ivwzdXRpQ8HomkXCeViqpJ3m2mvyHnN2
S/aNrXGh/I229Vv6Fei9lLmY22bvTe6MX+OOSmxJ3PrfF+PdATyIG2K7nwW9hGS0lasnNBiOXszl
vOKxkV/tJclSEIKon7NYVrKfPT4NKOVojj/5JJEjZ1cu+yoAdA2MpQ9/BHY65lm8tMwHk7RlQ3M8
d10/kNkeGkq8VK+ZURAqsllJtfmC79T27vnAWLc576QAnidoAyTaM+7SwgZsG49oDmoylGDw+V2y
SsadDlhEi90v8w13kKK/0AGB9LEgkWuql7k4BetF4RoWYRf85phiy8/GsXfxsDSZLdUJJUvPVv9p
NlAMtveROe8xHMfOco0mWR9DEWGW8ZCegky9rmkEVLDP7ig+ZMYMZAMjmdUsNjF5Qj+/PxbLYcER
jRFBpG9yyUtYMzLNJoKKljQwqERrBJ7JXQz8Uwtpxrze+cR5IslfxJAJ1qa8/gD7C5tDLYdLxV4y
f3VzLM6Vy4cqxTVZyAzerYkqVYLSVy0/22pRAY0++DUIWB1yOXQ/DgNn/Tam7h7p2hDYl6JUgAha
2sccMAFXVmF845uwFAktMKFYs+Mg79SKcF7edjUKkKcw46fi3tj5QODh8NCd2yQyfaqAWQFZ+kF9
vnA79RJsvAI2R1fBR5HTiAptGsdqn7QDW4/rPLpju5WKXLaYQhllmfA/Mp4lXc1iFKB+iM5a/qFw
1e6JFjzcKSSGr49/klVUvQ/ymjasaWFPXx9nei2FCeGIbc5kgCpSMU8SmnwQSE05ULLf6gZuOaDv
tc8Yp43F/lCkQOE+xzomTShHTV3lrOcJcnBDz+c63sk4Dew8EAbTI/mFls9XllFCQAKrZvjCc0rc
X1jXsVn67EbtLPkhpKAy2XuZAReYkrV4A+zD7WSbZvbmDjxDE4LdVrHBS0IWNv1lf1Xr2gUzW60I
h+jG3+3cFd2UsA5fobOO055W1SwX/FsXJgB1xV1IN6QCRjG4jnsS1QkwSUTw6K9oCFbc4zV16NR6
hWlRMueUonbYgUzo7Hp2EgnwBz+NKXMQ3HNrlMvwcW8gx6w8FTT1I9SJchar6tWg47kBlQ5ggKV3
uIcAGpsoErsRryoMptgTDdGlYlCfGY6T0p0JT928wEBSNadT3E8GvXBGrM8wFw+G8kktlgp1VLTT
aj/vwrMV8Kqxf0Uzjj/rL5EfkIetmYqpDlKou/Vw/iYgJpN7Nx+LXkEcLZV8zsFvvMvCn5pVEIfd
PqJZb82RW4koPRGqnpWRhB8lvZPuP0gXa/bRruyUB3pcD1B+zWd0WkT/6yjbggWgKwRiPJcHBePM
CfB2oK4egrORtWS3R/krUV7SykIWFwKMo96MFcsjLUedrNLO6np71FvKBE+w2xxYMlJIuAqnaz5g
o5miZFVgdk12aVVoBP0beAH0jTx/5y9SCi8wPIMJkK3upnurthZ159iTpjAiFrsgioWpNhg+Sj3d
XwBQkfEQW/EPPQWzCBEd4qAaqLscfzYAkpgiasccn4MDxrHyYJ8uq/KkKmtg/d5K4Y0NL7CRLmP0
4KJFoo1hephUGJtK2lY2MGvKzROgnYD9D0Rdy9L0oQB88fqdkilfoZzRSXKbHqn03M27fPydn6NU
KeSSBn/YQE4H6JuaOgYJmfyHl6eLejRjd8T4/3KYOGWl4Pc8eGFHemnhLtLLWhueSwsIBAkUL/L2
6FFCoyj1LvOtQ8RrNgxiC2I3a+T36SULeX4wGgmvbxz7SyfWANr/CkxMnXJRxMr0O/FQBHxCZemm
ShmG4BP5hxBYatmS9rX3s8kk3B7A6ASNRutr7Nc8C7PA8EhVUqu38G9zJ4HnnF8wm7i4YSujUjWt
POnPzv4flitYH1nQEbm6dMtEU3AeXs3xhr7ZFwcbZTIKW8xqwSexce9Tmgf0fy7zfYwIzY2uSsJG
2YXdIgS9X1fMwmDgOSpgzg0ggX8YqW9bzZb2cAjABXfVMtU7eGn+xXwq8K77GSHczd8g9AnCUHu2
AFtkLMmPlyrvrYgvcz9JuSYwTda4zbt0xRQGtxV5GaBA0rgMcQ6iHrNs+7AjKUUj2Z8HHBhV9eJv
USyDoOfps/zjzAQox3liv9Yyd+ORT+WSc92fP16QYy7/QhqLI+0457dfTbSjRENtk0tdc89WSpdb
9UIHnaQ3oJOXXE0i44W5AkosPgsjLDeVa7wwYXIl6tPbTvO7DAc1rHmyqZBRwMro4Xd64PcAvxoY
qUX29u8HimOURf8LSWr6sBKvjiOSTiQ6IEyIRnHLfAiWO8XrvwVezwwujdEUMLfb6k4yUPN77BgB
IntKkrGOwk6Wps+YUuYZhjtn1BEufoIFyrhmVe7AP82QWwJO8YMrK5V3Ufx3FtTW+8qcnHgxZ/Xc
eu+N1vYKoVS6B+XukXtGZIzl8Yfqhxidy2JlEMyCXmpEOHL6Hitsj0dGpVp/yfAZQm7DlLy/sbtS
L4v5XIdnT0TjtRqXuEMNZJxZ3TvC+AWtdiDUxV+k/gFfRpoS0QviPH0YUHH1SXT+tkeiq6Ky/gzE
+aoHbMjLAy6wqy7VXiBCqZhfXzh8KhAkTKq/Q0EkfB8WPhcyxPlGuk10g2oSjj46UYHgpKPeQ8/9
LBgXrhOXemRGxBFAyrJfzfItVhxPYbRLoTSG8/eAYc4sKhkXLqoCVgHdXHqBFE1TSHCUA4qQr0jo
GUuwhzQ9cwHtcWy6uMN6tOrvucOMQNl3NtveP30IhapqngXox86mzqSwwMmXu8AZhsk1TSGL9CyK
LMr72XvrCuia3jZtznSmE3GWY6mS3dsmggOpcJEtA8BCaLpFbIoSIF25YpvWh+8Gw1ym/yZ8Eski
qiSS6Q1kgZiBkx2yATVZBhM4lAdPwkTyRafehS7tz+D4b9yyn2et/yhZ7VvTbNPotSS98zUPEap9
wgEtDDE0jbV7iBbJVybgkTFx/ASGdoVU32N+f0fdzL+TbE6TaXF+w3lWiFDa3cI1h79B9a7XY0Vv
GZ/BnoC7TakiYe2U88GUcpv6hRbkgmBAq/VaD9spiSbpMglgPTit3afZELpgQ1FRZXnqqa3lYbay
oS+jZ2e2O+3NIKoaXHFOhgG2G4bSW2rFOr5JC3B8wDW9x4lafMbhvWyMBuDDap9dszdcSKiAIn9F
GUSrTpxYaIR22EGRe1DIwQKmUfjkJkmC+1E7h5bir971vG5gwA9eNfmDdTABw++P4Q0UfQlOPOqi
xtkczJM96wx9Ao4fknl56MrZeX9wI9yr8qK9igb70iurV8QihqF7jUXJGeMeLuW4pcfZOy60msq+
QcYJAYLIDuBXmIcttfEl5S+aLEnsdX/8X6wTm3t0tRfyLlffJOkkBtMYbPlCB8MB2xN3YWSx0EAO
sNfupJEcDAmkhZ/VBR62mqMxWFc2nPiFMHBoaRmiPBjDwtI+5ethd0aKeqCndgcSODeiFd0iQCsM
ysfOpFtWzGnqXTZJzsBr3ynHLTTf3ohXxme2tM7HXp+XUFJ7z7nQjauotWiOstcR/EQ12MNJ+l3f
G4HonloxGUSw/ShKHaBXvug5baw5lIpQIXz9uie1BjpIdkqhY0AHmAr9wd1Y/8T/wwv+BlagN5ZN
DuAKdLx+U3Dj2GmG0/+sn9YyuQFWgLwh3bQ9S6LdHROyTlBFEwJ77DIAYFAkFMfrVtfWcjoBDSAB
KMvUV+y1RloyzY89f+v6GnCOk5FVCCTerVhEpuESdmLcKko3EoZhGb+JH00JrN1orAhMLJLmudUr
4Y9/sdBKukeMHvAlirGEFnTOAJg12drvt7E+fydUZ2QKBgqVfaCDXLtsMuFexBtcOp0vFv+cnIKk
lDk1SsmGgpZKTm4kb6XwiDwKV8ZO5s6nraIFAzJtaLwJxNqeN41qHXRuyTyA7AoK7QpkwrpJq4JG
ZqCUYcKQFBabQjBBoztXludBJY2go1DbnRLz4SJBbKpRM5dM5Tuc5Vz3XMr9qcrB+6Wx6K07slbV
YwSR2msx2ceKpZEE+sLw9/0at+cgQ+37tjOPKA53lbAqUbvJTgAMmfZqQyGJzzIOyxX62YZqRSLq
El4TcZYB4kET6f31YsLXn4RZel8TnvPIh6IL0Y7DHZezsT4ZXqzFkxpofVGbLTb9ucswVpKMq7oS
pjo+qC48UvvbJBm88liasYvUIUYWM9aEOXpNGKenq3yr605i9xj+fdy+knKdibyZoV99SNobw9Wp
TGQD6pywpWMrKzIuZ2xK3x7zzkIeRyeTvwLlI8E8Mm82+o5Hwmwzo1sQZeUc2KmnC/zQPBRf3eS4
f4rtJ3f7wtjjZcIO0c5hKtSfbhEahGCooEPTqrskveTJGdi7KXTmxWneQgkB1RglHk7Z3Wpvl0ln
Nl1z6ZwWRLvNIvzDCn0NAWALE7b2Ra450N1Da1kvU3XSrbgAVu+yX6PDaPE7DCX8HhoF/7WtflJU
AzuHNlCf3SQKd5c3CqKoMTwL97dRtccy7Ng8CpstOwSuktCKnfHZq82jvjfGf/dwAcqV9ovGNve5
a4sLiIbR1oRuXm4OWJkXKV+Ya5hxIwscw6KqIgSadH3Ki12LorQ7AaOSlposHbLHer9bDTtF+Jhb
oF+P7eqfHUWx/AvFZSuwoib6n4dGumLngPfSathRGOTmATMoNgE9QuZwH5cR2de0a9OhRhD/4gZB
Xa1VcblLFCeiHE4YpoCNGRDmCqYAR1qWqpF+wJ0YkClJhNKXpGbRD84p0DxWOlT+vbc5Vw7FMHQM
oaNIOoWajq/Uy0Ub9GTtzbwv/W+XRytkDIaKzMeivPBMmRdgCoHaXOcUns9OhZT0aWRWkV/PYAKN
U8XRCrjSy/1ixY44/irbujIk6eILPBwWow3YQmjwKVWxX/JHAaoY/BKpgneyiI4qgnuTMqhsEVkp
1vmMIq3UuNrpz7g+7l88gIEPbHaFmocacfCHiMlmxsctfKKgkdbQWBlSFgzmZKCq4vi8vkPA0paP
B4XMJfOhGfdGLzCaWaaai4VoYO5QKFuXR0BV1jjQJJmcj6FUOwuD2iiqB/XkFefpQc4fGxpw60sT
Va6JuFpCK5hD5CcqCLey8DI8qTEtP2K5ALWU5d2UE3WnFcFIytWsI8HZ/o/dOTy6nE/oHh3X3NhK
FpC7ZUzY8auczXbfxiVYw22JQlEY/12r4FxcuiISaN3v7MiH4u3XDypuociskKeNp6HEEryxJpi3
zAgbhDWrIXflDAk2BG07P03k5VgUD05LZUCbxylO2lpzj0hBprS+8fuDYFwjsqXlE9NO8UxWOxn7
gVj25vbdRO+WZvNqtQ/IrT0JqsTTAiIUEFiXLrT1xHgOdYCyJKV0xmDMS0hmL0g1m9pPiAvPf9aJ
T06+wfl33xEPnQhy20HTFWizcwIlC0LsVsiILQzXB3m8+ZHQyFynMGgmwfWQ4aKn0Oa+b4elWqPq
nlmNnl54M/8U2e3a9SuwJnUkNjGQZneE3eNYzAkR5IB3opxEimQKZrUyIYl9kR6t/98ESc6zdXM9
CuQkTPJ+VqfjQJTawuSDRyDGxWXJr1i6F+8KpXgmlIbA9SswIR8ZkK5J9di3KDP6L7Wxhg0mqX3e
tFW8HuSt9PHQNPllGXxG86Wflu69aBsFN4fjmRAFDabcW6VRMq9BNkulct0LhA5AifObRIfSAeHi
irmd/CE6buu9JfF7DTHGMxF63HZGSUfb9Z+jNrOyMFtODbZar8zVAZI3u1jGWKTySeq/iD/gRIOX
dIiRw+MXI/Hc97RlYXgQ24Yn6psK83iRaz680TgHjo+JS2/hNtORl+SwDKzGlv5Doi4OUreBgT/h
UnGC/syGfft5RLxZi6f4eCwfiRecGJzcww5MuFyF9q1kyLeW//e2qB6X5erfCRCZgS2eSTRFqRzs
wX4sUjBF3WmoCRlZh9hZ6cB4vzcx/NtymGtTwSp7/aXPDky/MZQzGiqbxTH7EN4aBC1CWfrL08nA
D4O5nJBWDLfu/D4K29zyYytsmAsseXOOKxLC3dkGyFYWPYSB6OkS1DH4Q2i80WLiDbhnn+Tmmxtm
zE6B/cbzaZXaXAFoEUKG7837ott+z4kPxMtCc6F0X0doHmJPeOWMtQtmOLXhWh3YBBMQ9m4F6NyI
GXzbbfQPpdgbwaNcXrxUdh+y4dS2Zt2XOviuEPeBeu4gNCIaYaR5pAcieHY6NYJSJjLGR62u91oF
X1/MwU9mluPDppzDRdec2GIx9CI+plztnKnJCwbBEs8r8On5KYDBT5b4tUQSsgj1LfdgIGK+kPWk
cHjDLToKZh/aeSUImR4NBs3EQdS1NHpLTfdJ2ZH1g3nAmLo7+g87A0eeGwbow+sF/AhnogAUMz2V
qyVrppAiU7g24pNZLfnT7q5TINkzdxOZW8sm/n4eXIMLCvqhJ5VwFWTdO0r1JsKLtOHt++ZDVHau
eL564UNwrHAIyRKMt36pbQr4pEvvCX4m5qCeAysbHCgLIhMEdIXdp39Kg9i23jtxAgfm+j/01QfI
Ilo5D2W7hEFymhw5RZJnAEkVVd2YK+Fme4jYawSZTcnWBs/fs6ocEPdHA1y2WabAE2zqpSaF+Wcf
qtbAexexdsyKaRV5+PvImgf07hNZBGVhmmXxXoF9ICz8tu2sy/7mEPYkJPZ5Z9uP00VKAxsZz4AE
H6IZKmzRpVgrfg5hZ5J3y6AplXmRo/NV2mo+Jbzawfrz1qGBXNt/BASNix02jXBlngAmIts9jkAY
DksXxZo9h/hxOoW8uSFb0HixPta4VqL8IyyDrhx10E99hD6yY/tPvfsrNW0wURaETM5XFcomH5aK
CNtAudV57PIZixYGvBgYi0nPF0EQDlvjkq5NkNcqLWwnFXxqlXRV9HY2TZ7hkHPwt6CpjosZxDyC
iVpfdT1gt8CGvrc4bfcL4xkLpKi2vhfT9n3dQygjIfmBdRBxjPvb7wZ6iLKnAosPy8Y402OWgGKU
dFYFg6DREMZhJe2FoMcwR5riRA7YPcxflxzggHMcF+6Gjx8OWQonLT7K4ye0ATPOk5wHll2JAKg3
mCuVvUDIQoh31sOtZKJHunJckaJDQh5BdeOa6Mg7mgYchyhvwdSGvmDqXRN94HbL7LDEB1Qgqo5v
NzWnH6SOyBGCM4nKc+TwfUGYOVnwb4DbZFaar0nxdtzKGtHQRpnfw7DTb52PdU4h0mcf1789/vJh
lC7Ec4uBBI+L0ov5dUA60FciyG/freWP7xNfw7ERa6volRlpfILPJdBMf7t+TmRxJazolK6DvaUc
knQ6TCF6f3fUx8pSEY3WQwFD+nJkX5HZvj3+C8cqtoGjV6WoIfJyFoQMjMGZjmizpaw1gwBsaUrj
2U0oR/gzctRGkLLObchdrhFyYpXrLFRmVE09YGrQshZ0OdqBEPKNHjnr7mIX6Hrx/vdk9OLDIW/8
9Ao9N3KO2bGW70vqoWClmJq9Bgjl9aU1dcsJDbDiKzoHkONKGe+MYq4Pq0nO6h8Rz9+a+r79vo7m
46bkFuYERqoNTcGkIctv8DaggS68qysQl3+y2+BlbsyDAj4GAywPSDuYn5peiNURHrr26kABEp1O
ClHPGYRvaEf+bp8GfxYh2jxelss5n3qm5PAIjEQUDpEe056ldPRl4WP8kinIG7OGd1YydNJF19Xw
8f3tns/D8cH9ToR61b5g/8W2ZaQ9gJ0UXnTXQ/F0N12f7UVHwJ0kEYd7T7ZLNYOCMzel9MeZN1UR
/0X7WilEHCqLJqPosED79zuQc4Sr3gzRvQ3PG2HnGUrFbZ7WBLECbklYtM9qXq7vYv3zXPOEvQCL
LYtV1TaUfWk7zJioD/GGQuS6A2888Y1CLBq8su6xQAjO0IV0zMTn2Y1k3am6KDFN8ZcxpOVKpial
mTmzqOspMtFl/7aVKf8VlVyrDP8nuodWYmI9Xd4I8EWAqrUskVSKOEabl52PP/dO9/NuxUjVMBRf
gpoJHuDRk8JcWo9JPi7PxMAGtF0zMRwETyKxZq0XXfjLS4Te1lpsIWMS5krkOLqFLsF9NzH9oYil
Wkt35lyaO24qNO/IiRqg0e6MnqVs4w7ceQPFzNMOY8WAivqUN61Bx0ODk9UrVVXe14i2J3o/z5fE
z5PBK5RsDVXXOQ6hIRyz7Xx1uefI/9qCsZyQ4Tez/q0feORRyyiO+Ln+s/Fbw1lcgtcn0bM5oRhN
lMsCyzsPZJwrZ1ruXlTfBjkR1PuqeeKsjGeXR2UK0AyGmuq+4WWOJuKDBI6DCnd2K3oWo+MuHYPU
b2muqwufarqcmZ0gw7mlG5Xl40f0Qbhsa1rlW+d6+k7hFel8KSgjaYlu5Hule8lk8gj6kci4qo2z
QGaufQE/jQxNrqv7BQ4uGL+HFCt4jS6HooU/RHHCmeyITMFlAHqfGbr4rzbp++XzvNbQkhH7N4Gl
1l77AY7xiQRUrHwFQLUREn49Enbm0HwMMQp1iMMzDyczUpsIkCLhsFnsjJ96UzoPmzMNQEAUFfFe
0GoZMB1I/3lFub4YeAnJe6Vpi/KUPJte69wpYkaUVEw1aYIk2i2w5thek3zaKeBbvhl1x9skd66S
VMitrE1vjAagBO04zfu8VJtiv9lx8ESF6S+3i+XTes0MKksk8rD8DmvnTnJLfJ3RFtMsL44hsjfJ
A5pKuEpKp9yt7OBVgJ73lp+LvfJqaE3DI75OwO6TqDE16T64X0kCyGCZkSN9mBoZbijL1oZ2Tw62
8QD9SfCCkWeePPdidZgilDqEyETPXrLInF3GCh3iQyL28p6bFDJfELzPT5ve0ALrFREWGO6kRbS+
zeuCEn8pXjB0c8Y2ObviZMjvvdNoaFm4KRZbnppPf+jPXzeyMpRPGt7wI7H9E28k6RljYZuWIZjE
NpY/d135WRrENMXfLyKbff1vnuYKUFwQDQfhIru+5J/zYyl+211ni9Ho37QaRhLBktpf4Wr3KZ6x
KjB/EiTsz2QTq/1D88nPKNbEjuMnvZESWVrG1gnQNQkJDDlepkqJpEJwXV58xiYqQ5X3wAr6IHCH
4O1C4lluH1ecgIVQJmSAxdpRa+X6Z0nLpQFBKltMH7gZ+lwlbzzwOuohpfFXwCDbx70H2PJlYvtR
CMQSs8kc34V/w3P+hgGj+hvprjEBVRrhUWRvuSulQofrv880vFWNLyS1NAJqrq5U2gPT+EFDeWmV
5KhbvKHrgOJpiNHGjF/hlcVc7DbZ1/64zV74ETvWZv+oeOc6vIoAjaQxYecdXcxXAR0omRCxURVU
tpW25kCbLMf/w0+y7ctIstrRMq9HI5E01O/4lyXrtUL6VQ+wC4QGUu8czEzKHQNtBWzbl4mj32/c
QIef3LvFqdJ4BltLwyOHf77/yOhnlB0z398sxqft6S2ZKzVwEK9S2QFcH3mGigIJLhSE4bhn9wZT
aYXbWGo1j8YIak0YR5UUEBHYWxHonJAtDBC8l+bEhLZkqOA2kjpQtY5s/O+4akKIz6nP9Hg5aRtO
SLNWV5I1TyWCqm92uuY+1od/aLxlER1HifPx4JRJ3SoEyzxYvnpltFXy2R9u+LloibvhTSa4YOD7
LDQ7atSx9MuK3AXr0Ln+lDKEYY+/8cmQtWuN6SwAGfKCw3vZILIaXxdxLii9xc4V9xRcNrtu2fvW
yC0cUDp9JbVIXTvcXK8Rv6EQRcRPuhlpl7EngYZnwRIK7K41qtzLyuicCz1CAmOZAzpkuGcMKu3R
E1E5UsInzj30tO6Bg9MT24qz8fSve8KkJ08SA0FgpYXIrIjMgzWorLg7t/cuAql7BhzniDYawdk0
5GneI2mHwF99KtvcGGPTS12Yrg5IEi6vNt47sw+GSTfLMlLjYFGeMxh3gV6KkigDRvUFhUYlJh78
NesG9r3PSaG/COj03fSLIVlSleq5bd54S+rapPRd1HTu2mLzcbEuDvQ8kp1My7eJnPq+Q0/alLMN
HMxGEyWBryACiCTk2rLvymQVRKXoab49PrDKipwbJD7zW/6Rn5R5/whf5O54YuCmS/bubCUg7XYd
W1tSIn4qBfu/FicEicbl8iM9jrFuAxj7wJfZuV7Pjp6ATr+KLjrnAq+jrnviLxvSP9ITyd6+393D
pyo+ka8eZ38bkDcJOB2NYuwnTfNJU7a5/0Qoyey5rRIGjnhFwlXCSEsz6VOtWRN+0ZZzH4u0HA/b
60X05UIuDOzNteXuhR0WBCCy3p8ad2kxF0S76TMINDaNbU6eZcchvm56jFb3QKpDjjc1XiCnF5CV
bc18U80NWcz+OUXy0nG7eboEH5Ac7c322heq4cU3r3oWghWziFjEDqlyPZAzr0jQvqEXMTIVSwXS
OoaLvkT/zW0TnOE2nGnGOUqyx2pRthwsnRtL+MOcsber2MloXEWj3iYqq948RqLXTYZjz0FKlInc
xKVmMeEFe1IoeSpOcOlew0le77SV0S8NDVmtkB+j9KvDUKBMaNcwXMh8MlNggzJGmAb6DW1+LH22
OWWW9SxBNs4bbXnzfhWlzRjWsANW6q9dGWgcKAo7ACxBPTs1gjj3ALmwms2I/klN4unzoEsw/LXK
L8cHYflbg4BpP0rQABzBeV/ngAQrbB2VxD5sfzJF3LdCL6KpMH+gGdkZUCjLLXO9A8xbMwee6uxy
BoGwSxprTVR0wjWlHYquT+L2Eumr9DS7u/wY1OnDu3dQAufTNVRQLEmK8m20R6yTDxsXB6hClgEb
i2hQKYVlKGxpK1jp6HfrAAkg4x+/H1/s4KfMwKfo22/Dimk55qAK8LFricooJNgKCK2U9o2CYnlE
uYeBWIF3HJeOnLqFsRqVGi7/PmHkXBOP5uutzMWh5v/SwLL2Fayx3OH6/8SttV1sNpbNqgonN+WL
QGsMJeb5jTj29VwkEW00l/L8LmvHSiSKS9NJVDYGmfnFs0wrmXhB6rPAJUXGh4Deli2o+Mg9G2Js
7lRcLclk7XcAVlG0HK3FhbkHF2nRmoWDpLH3gkZ/mGauzTNToaoU6FeHprHtys8ILFem+igkDHeY
Zwf1tm2qZgWWLjL8HWlIJIUimHwuVCIkMgpPdauNgTPnAWQM2bckNhCtE/Cywekt0OjAqeP6TCxC
6cJLE0zUTZyzB+KEA5Ad+d5WoMU35J5NHZymAXhgDg2VFAAaXVwboYEOpW+Lp29LyaYQ6sRtYoWp
JiAMWavcr03mZZjuvfdmdeRxDqoZ3By9U0Gm1FIf+8oOee1uMR/vHyt+LZuZXym1h1c5GsSEmc9m
x22QkvYIxgSolCtSLB03MxLF73pZFGNZokI9vgZlTvHyxiBfFKkP5rjQOo+k4m4x18KItzru3Yi+
Lk+Ei1YuyjmS32nhyoM7+rKejNLRgikDbXyDWYH41zVEfaqX93KdtqMgXmWH6tqDGWptrO8gLp7T
NKlgjX2Pama3v7dn9T+zStQGVv25F2KBk38BKOpMaM5sIqcB/qUxlQ75l5Bvl+S9kVAumcFj2b0k
Qs7pF/bgB/oLfNnXpzRyHpsYW0PDjvTBJwTLqK9RBujUN4LO0uRyf4okIS1p+Hqu6oB06z/A3/hl
OASfL58taCniobA82j7lJ8UJ5kz50MDQ3w09v1H0P/gZVUBtsUynnmtqN3eRUIK6sR7kprljxfEl
K84R+bgZ4uKagG5SipM64mFOoLQo9RyPqp5JYPVgolVH5VAVRc/NrRvu8uUW6489hZe9Xx3ZrPT1
XpusC+lKquoz+2g0xyWJ2rQ1iLPS9JNroJp0lfOxY395b5oY3cRuOjvcYqlGC5N56HtpjHBFP2/1
l1tckBEWJujZ4TcO9kiuF4yQjbNpWzw9x4yOYwxFs+PrFGB8r4Hl+LRr1F7ZerLBIY/v53nf8ZjU
PcPvtz1UgwD4NISMm7TlcLl1HHINsPJqDVDvpEGAsquRmrsp8UHyDHigG09km5mUSL9qCWOBwX35
MonCeuNm+TPLgq+nBioT2KyIC3C+W5nP+rKyOLl261ZioCNwT3RiQrVWdlZn2Rv5jaYTA4YspUIN
V+URB86HNz9yNgssvVQYVuPg0EzeE+JLDzKrXUPxOzkrLiuSpwE2ID8YLtQcBWKq7C0QI/eToJia
9I7M0m8V1LBRWJaW6zEKJpS8jTKIhaLh31AiWmVc/MEhrsqyhhXwmTcOMKnspeKRkXX+tC3Ow6Ah
Vg+Z3R6cgJgPx2sjMMm6pM0PMmf3TR2W8qLbKai/Y4VY2+x5EZPGEqWnfhotSJcibZKmeKJKQcRU
rKydsY1U8Vgb6209jfN82MQ1UH2EUbqdt63MjHAIY4KbN90TJpEbtdz6AdZgNB1GmkFEyLhdX/Vv
P4Cq77EQ1O81tj+VaShADSk4EoLd/BiRUHOp/2+QTJJ/PwMyEuMRCmYgbILENIP12dPVa1ALN4FO
w3kwb4HjTZJKzY9f+m9jYf3373iTBmzoDcW/hdRIWaqUyxb3+IGzMcAP6Qf/FN/IlkWqVvDRNTBv
UaAarn6ft+IgJ6tYnXusV1vgX5nr/1VuQUWKrXnloJxg3sAshLjSc0h3oR02dxpcsHzqBvaKeowL
UE1oIDoGmL+FIlJuON8f4/jtFYgzsom8FUzH+TK61BPUsFzrBFHfDm0DTkIaHFpwPCdlBnGljzwM
SGB04r/w45ZnKjWVQE5Pw0XoWnsV8x6s8t6lLIxPmqCYp1mOzMv+K+CkCoFHGvdS3WHQyQ8Z2QTB
RgxOuBUQRPmogfAORjIGHajJ5+baPXfTxnNWK8e47VkvMn1dyHdsJW9O63rPnRwaIqdqLi7cCTgw
8M0B2F2NuCt9fFziWEUCtAK8C3/iGW+RNGgn4y/IBkbqB/nYwWSrjCn87vXwIclJWQTC0Fqe36+8
77qWR+OWV6+tAjsIAJCnQgWOsgqgkogG0W7cV225uTS+b2yMMuIuAfeQ8zPKS9Gc0MHCMM7M+ZAn
z5W8RaP7WIuSbJYco5lEwxXEH+Ld9GWwbqK/VSrKYUb2RagEfyBeITUyYA988re7QeLv9BzhV4g+
xLJZiyDa9OPLDANeajl6zYS+NI8OOKFRYdRQ3dbG07sYBYlaQppGPe4Om1q1mxPXQQkTLZAoAHsL
XAJzwWLF4Skv6frzTLw9E0h2kliz4GV+SvH2xvawwYOEaiLE3IEUckjY52v273rMT4MXIcqX+LEi
kLII/h029cdDCXZ3DCHlyx2m8Fu1t4wvVyrZ474PIJiWoBeFdKIVVNYap55aAoIPm18rXs7FY9qV
AEQ1eEnuzq5rdM1AzL8nv5/brkz4tFnhCbSTzkAj+ARkHYs492N5Aa5GKDTMoidl3TcDZv6im/vg
4s2Am8D7xWVLVtsQDeOSyZ0hGcxUkfcCokiABj36GyMVILBka16VzCMVVzIEJgEOyvF9eFEs9Vkh
x0eqnMEbAdk9vjLGbmkaw4HCtuJ8k73t7SFFtIDMQTgPWpQ6wNtNbl51dnJAdUyzQqdeRcSr21Bl
rrvWy0c7eCUgFff9rJ9xIgPdlMGLvgmbuvcEONs+dgGDXghXOmhGJq73VGi5uAZGxyIq5ABnyI+m
SGN0ZC0TMtB9XJHcZLVnPkrTqVTOZTBHZdJ/VamipN5IxsAUo28k78ddPXDXYgaJ0LXJblIGThhP
+RwU6QknDUH5q+7nEAYeTvUfxApf8nKcAo8CaPr3RZOlitAq0xShYvyMj0iMOoSR2kuV1FAm3+c/
q2MYSbVWZZxmkrUy8Jm2DyCIwV1tA3lS5lrW2qER9XFMUYrTQIvIs+RLDr73KDfo284GVm3DYGw5
exrCSdG20LMPMgP143mIR8Nbzib0pa1XU94A+M/vWF3m+XABYpRBZKT3zVtcFUV0wreSSDHAGua8
NFZuGbq24I3f7xUL4TTIHZ3SdGooIBv0jY08TCfNCcXAEvCBz9TvWrq3WLHeMx9kACGjHR1vzqHe
HuEtYNSg4B78A16f4q2oL1fjkPrxLw2zMoMQdxReIfBxyp/0dO3ZXnug0QHogbxvX1RgI2Oj4+f+
/z9zPb0rKe4Krr1lQcS38SBfYRTzQ1VZfp2+f5D5fYpg7zgufPFJRsdT+nnQyIeTXojFDlE3m1jz
40VOVrmi8AQy9wuXR57zEkHd0cIvAgAwzMZPommBpUU/zT0S/mdkvR403orTnUvG/VNgubF3KzrV
NdKqFt+LrENI2QS1bKorEnnhRfJ/oCxwYQUdecfC09R7T13B0Ru7dqeVHxynS6fEk/kTAzs+Hl5u
ASp05vHY+oVVBmcbtflYYNOqSxefbaeRrwjH4FyuDaaJQ9AUWVUFhlsh11XT84XDi91I/Nax3xxY
F9mxwzs5E9dikyb/5Ag5nxSY340jss8esOKd8XBGLHOpgwcdEQ9bY3IU4Ty+sBiyiOfwH8zMEmB1
Mhi1IY/n3HThQ/Zc55IuUOW+jga4hRFRDSjxZQZNMK8SLBNMk3OD/XipYfx4rjxE4jkYqM2WQF40
JnsomZdy+uoyBJFaZwcO0FmVfhZ6iHZDVWFmRMa/gJm1kJ+rSazCFuhjkJ1Ww+s9A49Og/QPXn4S
gE01I0RfVLUpKjTPSmT2nV52O/p8br9z9qPrsaMy4hJMOrwVIMK3vs0/rHr4tc//soUsi24Y4kWH
kO84I6/s0RHuNjJNhAzfwcxaDmSdKy4A6LBng/Uy3oH/EXAJTaRiDFCA0T0w8fV5gOj8/9Fyka29
03ZNoYxKM3cuLF6c1/1pPx9AQumd9fpUeM7RcfROZTKxcqI6jKEM2PnntXgZ8BquIGzVfEsXn4up
ARTPlC7icvg5JoXNrZkfdIyTXMmoCfmkpARkt/q4xvRyUy138mHzP9c40pU3vmO8iO3s8AAe1uAy
ijWaQNywlkMENWMhqqI8vGaDnF5KqQxUdgRr0GvWWl+YAfXUxf8y1YwPeLRvcqBvWqsdG9zU7j+G
iFI73z/RbQ16Jvf0sADDJIXEpH9oU2KN6MRCCnH8b1taHxHiSZ2S2a4cReF7EzhLUYZuD/VuZAUK
z7An0HHD8dsix21G4ePGaCcB8caTq1tlYVnmWiQ2t1eUmsyxmLOSJM22YMsFGfQaDv+d09LemNIJ
zUEFtOIhktK9ldsR0pgwcPLzNsR5IJZJA0+2t784rz8KvNTHWpQO2o5uO5XyN0ddoIPNGC8NrIqO
42Xe3pZ+dcDkoroBd+lUGZxahyu+dGPo1otcaqfYmXHQiGJtmUVR2eNIVKKcye4uCbBc+JyeSw64
PbCXyid/VEXrGxpuPYiY/ZenGmffCYst9OMW2VuCGQbsf7UCIvyKlFV8sM3PdTNAPcoMsAJKYzRd
WQTcClE5Uh3UNX7Z2aIy/YX11hO0eOGi53ff8c4J21ZNh7vf4YXjx9E5tF/opAeKJhivvmQ0rlYW
/+Jg6pmC0jcer6c56XZaUftTc/oCLRItxByIKr2Uh9sJbVYwfRme8ahv8IId3f+a2iGTWg9Zdn0x
ExdMALUSaWEzb/fTXMtpGpheD/f/Gpa8mJrLjj94u8swYp7dgrjeMgw5itGslrIg1owu/7n5wDZK
LeZ6FzYGHgEUbIBlWrLbRbPpFwkDo9A+9DQNTGvdJ62phzJoNy8z/O3z9iFsV9BymGa4NLghjgdR
pAOdZR/ke9V1m40A+EOFTngXBl8XWf2+b8LyGVPvbhlE/GD87GoUX+2JwgoPidf+686/j4vNZrJv
yz8rbvznYUitFz1K27mx2utjvOkyF9HSsWJS0eMPLivfLUQQlolYHenrAfyvzYNPNBHcLJmg9pcG
WGhWUhTiiMVgfOjjenpHO7nCAy31p494Fvf5e9dSB5FnFwOegyZbFKPiRrvU6j7XG10K28XEmWzQ
nKh3CFzhuZ7Hjz3AGj8YhmFZinA2zk59kCl2japjckXtuytMAC0L3G28DOYaQNmln/m1K94sUTuQ
YWwB2rgecM14sKc8qZR3B1lzr2oPOqvzlM4xR4GBVWv2+ymvh6mKmjBNBAlsfTHdSJAmBlX8DYbi
0IVFfSKpGnDX0arto7q9Xz4Va2Nj+hRsSuGhrdxo/kica2CgR4MiFey16FCBhrCMVCE8Q89lVFA1
ijPkqOn8bWlUi/Z//YHHhaiMeg+7gwECzlLV1wQxpQsJl8ECQ1cvL2V+BOF8O7+PUlFhzFXOYH5H
13uiw6kMfy3/mlOM1KJOZsgbgAW5ltyJ4X7p85z3lsPxtNzjR2mlgCvVKxZXHBBDVr7YIYPGbyVv
pVSh5ISfSMRHZd/MOhiaGkHcoXhKlbc+mUIePzqmOjK78PvvEmIpscF+QeY/u//bD8z+21DFTMwE
tVqfm7nWwPkPf9JQnRZw3QcRjYm44gYhF+pBJ58uOQrmYzVJaFhiYIXkmbFWEEG+vBqo5IZ7CjV9
9UFZhd9V72/sw69zGrs1Zca+xnTVyXRRn5woGlu/jBM1oH/koOs/BXSSELMrmGKp4Iq+J0Z9WvQo
+y8/ZraQvH4e5UqYpUbchlpIWQ5TLm0ZLNwBGJQ0MPMJv0i9hJv+y4GI07CFSLHhNaHLk8XmxJDN
Of8pGF/HrnxMMA76mNZc+SBVYjrDekotz52EgcOUXSGdLF0SjXrjdakzFGBJlj5WUVgGPSxCy0KJ
AsPvah/ck9xIkCqdmiYZAU7xnHYEgFTsf8fsiVv8ds11W6+p5MdOML3f/SathoAlxwggJzSQMfYT
Bg4EbQrsPGgLLQZSZxSxnDHygLM8bVoKK8//KyPU8tKUL3xtkl71gK8ot2TcmKVLypVFNcrSjKJP
vn5BYhHZWGvGoxLLIOTO8wS1DAJX2EtqhSccIoGRcz1MFCP6Fj2quZVFX/vnvaEFSObQ26E/c8nR
2+sbma8TICgrrUVDt2UFpHbkVY8s0IYgQnSdxNTzo3pyRY92iWtbiwJ5T0TjQwAQSHrnnLFsJWji
bLQUFi+kp49ncHMQAQ/4gkjZyhNCgIOhudNUO+4ffhJk5PaIGLOqY1by/6fLSQka5XqmJNMEAGog
u0+VPv4iURilzJTMHhXjiiSy4cSKZu1luZEDY7JFhYuV/clzTIqQB0eKrZF0GgyyMLqAeJpH04WT
NNM8f9GbUQEJowkfNalA9cVTjBDBR+fLYW3PjeFx43OMCbEdcxeJZ+yITA+6ERSOPFzinvFoB9ki
zdVJrxKk+2QMLSYM3AleR6xn3e65yryZqfc804tG8F6uxxyoOfBaLybQQaEtqB8NujeGTWa+Gg5Y
aiqOBW3vAoKcNtKx3lp9en4oHSwc+SjZryHP6UW1ES0QsoPnKBBzEzght190QWY+K5UaFV7/gJ5C
k293JG8lBRW7/9zqiVF3DTtwajCDTuDLV8eVTbk2l7HeAU7GAA3oXWhkNPiM4+eErA24vZIVbkDN
ERmtyj6eBOABuqsYOlCtueRbOFJpwDhaLh/4MfwHu2fU4yfoOZbmaiqwGbmhJwS6zPomiaTKB8Bi
1viDIh/ONZA8uMWqMEL2Xt89OBL9nukb1d0ohuB8bC6ztFJe4mr8cSUPRKN4evs+6VAhfOBh0uuS
Tt79DvhpGFlcFM8rsNrtS668ADdZblpb84mEuzwBCxYzErVZH5UQAvJI4VvRt3SU77SAkG09rfaw
JF9i/2rzM1IjsAiiewDi22JtBbe0jxJllJmH1VMCd3E2GbYm1uRWrUmqES9hunsIhosH4QmGMorC
CUYF3SApE5dAGOpHQGegzb2iyj7h+lqN8bY8TMfT45NHv1VIIC9va9bMuXsVSN5AIcrQ5AbB74yi
YB41xJ2a6BZBYgsslciEiS52lbv+mgXODsInX6jRV8TkdA55yAyEJa7A3Mu/c1U3bUHqG6RQoSVb
c/rmhURa6kPgWt3CbjmMYLaRHC3NAQCpq6I+aSU1xbUUVEJCDPUYMEBary3Gp7lSJvJmtWOkKjSy
XoOXWcODY2thpSqNfKrRJwV4GOpYKLSzKe3n6QBiEiBEhmlLQMCvZMl0ks/W5H1IzsWrHb/IeOSk
YRLqTfXZKP4zBykYWDGFywkfudCw0CnYVt6SVg9lQa7TzTcrESPSkXrhRJqjuj4GQJx1WplbKHYj
N3nHrfmtoEXiQi1cqv32E3PX2qgH2Albivd4P8I9mjrBDNUkooqANbp5yBAQQwwi/9u6REpA8/Xq
THS7/6HjbA4/xnB9wHgo2IvOtu5OGpswE/MduepMHodq1Z/SPAU/MImz81/4eiT2ddJBtdbpww1D
Ps6Y+JPjnRKD32RyFrXdpjL5mDsnfrLAhY+ter63cr0YAPnHKiFNsIQmESOsGSuWeMpZOysbxozZ
Az+5qx9wwesvnkDcu6LYoXyEjGp0e825pMZ0TDcAhQL8Jb5gS7ZFBWR+779Ov94Yzn/fOiC72CkT
u9S8QLMTMQpPqFbL16pcoYZtzo8eIY+2NBzK9rB8jhtDUfcqDmxCoBRnv4QXCRfJiRJKWsDwgQpD
mpIGosdssvH4ppfyYJ9NF6G9IZfoU1dYOWM+X8znVJuikZDutenMuDXxiwiaaFGCrc/9t2iJHYav
KfI4LOc9FFVrOeOJD5179f+BOAjmSpCCNO1Yt7a7FjT9/BtQCwylsL7KLrdNuvzNYwi1kh4ykSLT
CAUeZYa3N4UzIsvvNe7rekWVve8cH+5L7zUIYGvuJF+/o/+XZpIJAwJ0bB0waQMzJgdN2+FYsQ47
HmGZ0/0fpTglQVFNvcxMTRpueerODYJqDhjAenrJ8v0dXuRdAHBVF07Y/x3XSHm1mS+vMY5RjLf5
5iRtC/vPAO6kU1uZW3HoItxKoc/1SPxrOQ7sfX3Bm/q1atRH6CMM/4MpOzmIYXL6awlfQPqsRjMs
JnUNHMPoyKJmdXC5s+PqN3Vee5v50oH3P6j4L4u7Af8dAw/i2z/tM9w0vjY2OAFtU3+xau/JOdRm
z+2xiGaajDVvAQnlsjosV+5vvAcqFEleyAGg1S13FhVUCvY4ibDFH7MRWqv80wWc1ff8mjLw5618
TlhZd+YE5IMSt0i6YbWRjV4zMea+UJe5ktO2YApku5e0MLC+hiSQ80A77sBiTTDmhXv0zq/0G0nc
bLwc80zTfe5AH2TrWvVqaQvAf0MroM3kfBwSfgIrEqKGxKkJcRbbnQUORlkQ8XVFV0qCPhew/18u
s+RBtO1OHto3ztfAHfl1nc/BvTxPOQHfVkn8JLsMoHVsZ3Xdelw6Bb9Yqm2muTFHOXO8AZRWsyRK
p6ta7GmeckYm+3IucNtiLRvbG1jE0ce39NV7yBxtkEodJZAqIxlePOrDwozCU+ugin0bIzwZ8usG
JTKdv79V5QW5moRRHL5zYp3W8e3VKkD82SLona8RDyNjZWvnufw6E8+7Idaz99lA+7tkZWJAF1+5
bLsjHWdTcXhAaUGMsNJCCOo3XqSpGsbi5t0r7e9R5Q1oPsBVu/K9lwWSWnYGFbYcPldsPQir2lPO
qpab0yi2vaHgc0m6OF6lj7WnP3ZLvZYig41gcYjiVIfjyvWrIDIMXCLsDeXvNehWdIXAoryr4iAi
KU+kpRaAwZ8S0HtBCaO426G/mXK2Q5Z2dnRp3fOfwz9pzRm+ovp6KVCDHEFHoBAFhFI1CAdPBjjC
BXtj8MQgAVk93yZG1sM/1jsy1xYMuD+dbSudEEc385BbZuHUKpbRZ407LU+HD3oSyzfr9VCrkeG5
GofuH4wVVWEvlfJdAI1OaJb4MuG4QDSWbkgWSjtD1X4ZkG1TW6F+SrjJSSsnhnknos0CsqguMGJ2
RZtg04UbHN0twCNJYIlmBN1227XHse/6MflTjTgg+CMyy5zkMRqn/oP/Bz10cJ7XQ+jlt7RGAwkb
wCweOMofMfp8yClRmGIftb225OEG23qBNo3QDlSPaj7PO19GQuXmQA0pfSDtr6w4AK/7BGx5exz2
JTWAVxQ8DfBwxAKh+I+JTE4JnyWDq3sCtzhJ/ShfIqr23A3TzbtutcgmY/cFP5/ja78C3oRpI3eR
6XWDt/Im3YSyM0vHW78acmFYPtfvTq2XAQNevLjU5D26DVc3c08j7E8AYKtxE8JpirtNqRPfU29v
VM/wGq4Z54HIrGhPPrwLLVgtFIhhrWuTVJRq1rzo3gCMiGSFmDA1gUA0AlshvGHY6ie8Sw43cdum
wn2eGrDpjLq+WexMQR5RYkAmpoNONgMm10zrsLs2FXHOuNhXdMuAzN1zLeG+gjWIGTI5awOag4Fv
Er8GivXoC1B0c3i+/OX2opLa+M7FVRNzY7LzHB+AnR238BsILKTFJV/8e+6tk9iB1KCf/J1GX8X5
bNHEbnZQr1BTBymcFARd3cK4ZnBYpCgbFzHfvHb0AOvDgoPHfwge/ynYQGHsG0yAyNLcGt86TF7a
Yzi2Gl68w9NTROw+5fOWR6Ajn6z1PrwdPQdjNzheYWSmEblXaCr+7GU8Wm7R9K7kWcxS73CDi8v4
ymBGSA1BhzXnS7yPihUORCeXUsPyNIrsN90O6njtxAm7CGG1FnkQpuFz2skgvcCoXiUBw4NJMEf0
vOLsvNAt6S8TvTc3xNwFrBW7S5xGBBhWXmLJG9BWFcccfOtuJCU3rtAHNngBzOKLfGPDnSk2riV2
2bCS4EzdefmnUgYZuo7j66goTVERcswk1gLIME5UT/+0YTwB32WA9akf73KogRBg9m04cYHnUefG
M1UoQoGNkvvoku1P73lRchdgY05CKi6tLaXWV1Z+3n4+26SpL3nB7/yLfyWmpnMvrLrPOpm5CUph
+AIpk98ZBCSvwQIFarpxUOgSmT+vH9WO6FfZhgmP75ohzl985MHlTqlBnvkM+9eU+8IGOAEN0xp+
oQuxOtBwNcUQpS0bNa5ghbZo3fWSpS0SyvewzzwTK7IrFw+RyrRVxBl8pWzmegUml7th/AWErlPu
q/Eb/Cu9XOIDBszawqDAJmrnFmjHVXGIaLjwjooLV9S5M+eLPxwYP64Pn3f97rqprtAqN37rf844
o2uH3pbjP8x9jcirNDTgqobMHIRT3ipWB0cP/vPBzAu7d5KcDk+DhhiGsTqofx6fdVKsoZn159CR
UEgIub7kIku4DsWPALZGSwb2KeKQJrzUYdRwN8muoUPeQzHsHh/ldpw46NleyIHRuV6l/Va1af9l
Rywq+oksMJ4geWSeynuxqKiKm77MAsQOPWNo356SdUGDhpJIOamOi6W6LPeHvwCKNcg3RSkT2k1c
DLtaZK3Nt2ZA9Dj1w1kYpEYsPSbTXV1UTaeBFk+KJG8m6xocNcdXSg2YsuR6zIHRR8gKuyPBtdrN
uc4IW3mXfEEM6/olxXF4XzK01W5LxzcNc9dPixJlPJmmNBzj7DVfiVyTnzeg8Ena7QgeZFeXUVQp
50T3N4nAlBbD2ZG/y32gegZOGCHGj5SSYTW5y3oXWQCCrwp19ME7rYh1yxSjQUsDeM/EhXxERBDS
bmSawcr0+JmuR9+I36hnvicx2YHyilIa39EWWVSf95EtNFsSbZQ13dkpqi7C8s2/30VRp4tEC3E4
+hchxuyz+8F0xoE98M9R082nG64xsnTL/vzVvytYhrYdtFaZKAeCvBS+CSvR9Yj0d7dTBEOByttI
jSjCnxjNRqtQV9Xd6nt7YZrXXye+816ehvEyQVCpM8P38WAZixd9/7nlvR5O/z+GozEpt2/dHHea
7aK/0NmBFvIUe8lwUEqRv3QBlivLhSkkD4T4vqZO55luR0D00S7exbjxKcCiXOleGviHyyS75rMH
VMvESX/17kv6IO7Mde9Lc4uJcrEYdamxnt66e8rZzszCsgIhd9yXT58tzuuncq4Kk1818MJkGY5u
WqBNa9wffsQ3Fn626Myo3Jalm/MHzaD7r27oaAvOI5pv/iYdq8m/fB6Bfl1cfAY/NJ6O+X+UMqkY
+DlfQIA+dFQmCklPBLgX9d66bWto/zuE0PEjMt3dV0a1NBhDFDlchbIS+86JBqjLG0+MTks+rWYa
G/KOy9AtuFDi39gCHLgDDpCZyJdVSuIqJIl65vEWf879uayY8cxBtxLIlUicU8I934QmXnesRH5A
cXTwMRHFUccP5Wex3PHiHo5ebOIe+QQvtdv3do8mYR7uDk9UY3Xccaw7iXthTnO27R5Fj/9gFGh/
5Z/Vyoh8oNDg7+GG7S/Q235hx3HdM5iPDaMcXo5RF4b1q+1LypRccb0uuK937uZuhI41ks7Hk+AO
ZlJbckPkDJLIbo6D5RnFfzLHUivQDwIrbZg42fxa5vPREqWiObV9lFj4rDD2nhYyssXabbpgIDmu
s9xbwX72Q1OkvlIhQB4jRv6MvaTcsQC/aJ2lVELegarOcYfU6febzeGn2bbAKG9/UdeEztxsoeiL
zqXzf29kZQb+Bg0BAqzMVAkajpDpJcES1b9KUcp/KN3/mDPTZGTthPbJPCwLOfrH+2FYG9Qwrq13
uun1tnl/W58I7Bnw7T/dVDMCXKTzJT3xlOZNsXuJgyIKhf0PyuBgJKX4gwpkEHBFbY9Xv/4oprE0
DA0w2WbOeeCK71PqiqIYhOW50X/3qXJks11Q4oE8GcBOnKx+vnjS2q1wsOx6YZLQ0b6R3nS/a0mF
AYcUzg71e0MIoQPALh0lhVkTv15AhEbvDthF1Zv479kDxmG3XIEOUCcBvRzfUuyTgolH86FCxc3b
fnOjpWIAqdx7nBSrjJqqjvuJmEi9dPd9kWpAuz/jHpTO5EkqYeLfB9nqLtNWITZrJx0VFkpwFaVx
MrjQ8GTWdY0YSoq9yRvOkpRMgNxS1Uy4lRMpFxM0aOohLEfosyspINVRmxRRAJOH2uTlv63uSqB0
y0BEAW+R6SkmKJ4tV9zJe8yxL3CeUj5+8FQXUUGCZWXsdzik04c7rvWwXGSPWfIBaRQkCv38pGej
aXuPiZGV0TTUTVJ/wW6cmafg3kb3XDf5Zuw4dNN6rVsVVM0lhymVhOD6agTk3jpo3d/0lAcuPvQH
mJO1j43MCRV2mN6uPKCgof1hQvvB2OUecwzjws4sKO40HcT24Juk0O+DCUNTfK9xoXr5bC1KDptp
7legP4dCZob+3EVVeECQZ4xmJWzRuMytXv4dAH4kMHM9fInpA06GZD3O/oyVHG0qP3NbSZ2HZ3aF
4/RmD5VTwKe0Bv56qZWbU6dESnr1jt6qXpznnNi+3sfa0SRocezF/6MCk50WqUmpQkuzWO72VQTT
RZ21xqbiI8q52p5tq2fA0Hf2iDdU3KUwmXzBtxQdeF6BE+gFofTgU514Xrel8UDBNcOoAapTGNGX
mSlwyJHdCuGUgpYzknWL5Cq4fslv2mhIHMUScXEAi+sq9tsvPj7Sw/Epg3aMDIG9vi/t8Ygl/xId
Vq3jP9oD1+S1zpxrzXX2T1EEkzcnnltCE4Wz3BBpXCbwMIJY7/sy84ko7MPLpghIwRD0HLrEuQEi
PniWWGPIaf7HGgA4TwDa9jNq9FRBWGmDe5aNy7rActiQogSDUfh8mSmgt73q7F/6cUw1Qqxo/T3w
qJtZepDCSkSNAE/5Qqz3XJLhC4659kHv676mc5RWdrBix8xZi4L2RkEJjzf5ckJTkqkOD8s/LU1/
CmnoNxKzEwy4MmsiCm8axmtY3I9G29YDEQXg9oZ/YWWN2i+Y6GBXlyzKzRvbEOg/o5m+FxxBRJRt
Eeru8qcWFjlviBpWtaQWrK8mhUTdXIVS7EzsZVGT/dJjsOuo1DnNuYE6h3f9hlCNXwJCE3M7Knkx
d4OcgPoXOoRmkC/HDWoSdtvK8JHPS/5yyJzazvZ2myuX2KRZl6vdu+bvBs0dxjBJRbU9b8W7kE5g
xH/3IHLXwVMrFWaG3rvV1JkuBc4/2TxQTebpIe8Mv7Azh+h1QuFCzXgoTthtWqbbm3tVzSeZrGaT
p797XpwJFaSRWQHxAU3dHI0LHg60lN5kAGpbHbDHJrd6JOP2lk+R4NrEj/Vp41s2wiJENgzUymE0
cSaKUc02Etro2zX7gy3iz6/Lidn7NSLFgAoagYhKKPhQ6kzFnaz7XPFaIA1xI1dP15AnPO37FAJo
bIHLnNalrd6lCXLgLMzLV9z3nOlw14MCW8YJ5cfd/lb7X/+XH78KU2SQLNiNUp6bfI5djCXp1rHS
X2k5rc/C8flw1nGaXwhjvZbeAsq3tBFGYVdiFw9elV6xSX0OSBry1zcdoG+aIm7rcep9pXdYr+KB
5weeon3Icsq2bhh1cOTMnxFZO0tirXaJczKHnM76wQ++JlI6qGZ2hDznrBNh5YkUPe+bQg5r9XaR
vAV+twzNskvUctrsyREFugj352nSVoad8BXhBWeU0emD3rEgoSa3SgDL6TlUKkhcsDKrHS70cJyI
XNDmTFxu5QIvi+73nzou1ywqGfh6YBA06X5vDAG2aKj/KLwBjKhfsCz/xw1KDyyK08k6ZLDrPrNv
W+O+EzFuHaHfi19SUKwj1wdoYLMYNzKjI+Hqnd6fyel1KrXZk3balM1QUm0EuKHn6A7MQUP/fGL0
YUMXCyBXUEmodkoIBeNbvY3g/cn5r7+eq0HF+UlcaT4DMklEr3C6gCQHRCYU2lCL93t06EGc5tq7
suM/mo2A7gMMrW9BmjpeIT93DD1vqJ/78z2ihiF6teT0BrTkwYn0vZtqUpBN2/ffUNDt8Xysvn4z
Xx6E5bzV/M+UVM71tY2wWd4OEQ2hh66eHX//sbrelGPFQLti8srfWVSLwC9hw8ZZtJEfDap3meFy
ZNn2egV/WQ1jXjvPwm6Emg5dJKTo28KMxgZ//mBf54XMUNb+rsJCT3n43cMxdsrjemA/aYRF26gD
IbO+cBRX577Oz5YIXj5zqNxMK76n5uM0AcPx7nQCyKf5lculDVZafr18Z6Cp0qB+O6+e+jPFfnt6
7pvgy0eLVfBxQYTDfv7LdjZQdq7zuQCi9OC5Mv8WgzIMLfTXZ0W/U/IoiDPUoegVcXcv8/JaHE4O
vDPx7d8GRVIB2/S3Vk1shpkhEijYgLYZemILRMVqlud7meVqErrhMyFiWigTxOOz9DhKIf5lCUUS
XCWRLGikmRm3h+Wj4XzMReSgGa6rIghZONjckJExzmlXg27qnuiXJu8nFwLh+u/5fYII2pGJdlFK
FJt1mSTlOtnqcarnqBTTv7jnX21Tk68+TdWv5epEEXXDxBcY+3kgHM2xkh700ABok3iwHQrdCJYo
Mz+A+yQ2wAXhW4xeG6LLsQbK00z+JwP9BeydRImL85WXR3AcalffuFxhRumkzKF4qlpuapw4iGEK
Jzn/uykiNrA/VEvr5X/WYiZ3XLYVXsCA72CRdRvVKRCoVohD2VsDrUOgRXd9A/zdeWEIEchPC749
slozkT4ZOxxfa0P2Qz1NKb8gtvv4MD+/Srg/h3UsXat7yz9KnSHkMdha8B8wswW+nIt7gWP9h22F
9z4UX6hy64g9QWawI2fe94FEtZmWW61EHzCLzYJDo4/YrkSaJ/FvWvx/yuNg+n61dN9bTamscShA
Ce+7A0g2Y5/qV5C0wAVmxkbAuxh91Kzp+NRBFvXuoRgcIDNGSQHU0BOx4CoaMf4SckpNHnK9m/ed
RBW9QIuULSJprArNk4tfC1x8uFwvPU4lI5YHMO0yo7/f5MCD1l2vvVF0npGNmt5W2lbSZf+XwBgB
+G+UOnuRBGksUcRhCQ1wTHPn7l25m6uvuSF+Flnh3We3EbJSDvhVd3Rw4uAzJT5XfN5aZ9nFX/9s
upGokx3RkfyAwnoR7S36rVSBFbbosbvKNBqd6ZquHge3PUPhw195wOyNRqwX+YelTZa+rSgtCgoY
wo+kP0yc+0xAqyx9XXbX/SjcA8LiuXhjCnEz0M4UgpPIyP7XlQ3m9WjPbNhqw7N0Mo/MUUFnV9YP
8eOyDLAxZiW+UVvvlJp8PKEP/RJLMwQ8ZCZV5bIsZJEZlFmbcqCpy74HEURz6PTOOrWRnKKPlDgZ
zk+Tj9OWRS0bvRJJgNseFd/OGyRIqohHF+3UNJeeUy0hknrvaomsoh/n2cfjWWK0HCvgslnA9tmC
vv47wFaC43edJJfyoaGM6RaZsLUgWgcvH3S3nmx4+KxbdCDioMIt/LWcx4WJJVGyKPtykAvP+qKu
RySj6YvXi7UpZCuiYYFZ77S/WM5Gk263pjdEp+Q4vaDS3QGQ3H2hfF13T4UDDRRojIQU+ysmozVS
kbiAw65KOEEL/LJds2goqH54mOJenr2xEag5+UevwzlCTlMluI28GjZ/lRfagLE+AOGDDyLiZgwA
dthj89g44k3jGnYi19el50/ekQb7tlfo+3siyf6ttkfq4kUMBgkoQQC+/mFYHVroOFbugd9L7ZH0
gh3HQDcD0ETbalToH1T0OQ9pZpv9XJuggq3Z70OPlM5zPPJsHa/u2wzMEqknzzSMWGzhIhSlpOq1
X3zOLakzLzgno8O8hwhZi81xmx2a31EpU+M9e/4TM7Bh8xyR4tH6YjoUr1cBGT+/rWzOknp3LfV7
dBBD6IrTUqghgsEqF4pY0HxKEc0Q88DmHz826ATNQVXXREtKbfGO/Ekwlg3oHKcQNkx+bYJrMfVZ
9e4qZEjfGaGulUeTdB4YdsoE1ZAvh+stTBTvzp9yk7c9FG0PAYWKWoxzrmZMCgRK2nryBeqTtjF5
dFErEDxNDb/CbwMG6g9QU85T1uPFb0JB48BBhWK0kUmIs/lIheV3PlOk7eGb3HE1wiL9PSuHKPn7
jQecK7nl5mALlYhxBfzNLYpWjzsb7KnHGZF2cROMVs9JSu3PM+3+AY9OBAlpiRPZMPC9/UwyZabu
na1/FrFnls81ueiUXwWT92LZ1sVe3nmEtCsyXzUxRr61oFYCQLSfWZ2skuYbyh2/Eiycd7AjPteG
Mfbj7AKzSqbX3TiluAcOWcopIRuQ/W54tLp3zwa3tmNGZme+BnrMDafxNRQOe7k/NmLMMSIeNnFo
nVH1sUUlHQIe4c3bxc+T5R/oo0malEkrzi1TSmoBGvqJKuc6BXZAbVMPXZEVNCAMMgN2xgMuAXQK
EHhnEeYlSooJBKJ7T9wRgtZ1JZ2tv3n5iPbwpik/cYnx/CuiT1HLgkwfzvYhXjaQv9VBdVZkV/yQ
xV0NxYHEswlQEKrDGXEfFel0gad8kEQZfydGOMyNblyaT+Ka40UP96hV0JgFqVuIdTY5ljrHe4ll
UOPbfoBKL0pSqSvtHalaKuFrnn01+oNS5F2XF9w6MJIdYWPi3xC9+OIoIkqCNGfij4hIVtqHbMuG
/Gmkj0fW6Chc25+RNHM3m5swZ6oq1lRxne1CwH4pmqubBcCZ1iP9XFc9+8GljHSe3EnKvI9PEWes
E4rhZkB1bowqOuA2+EhAhB5gGpUmJ11WG49HcRVDPQAgtubU+JR1fuWzDkdLgni+/u1MMkf8ph+U
8W3u8zaN3yrA3/0tAz8S/O3kLQlJVr1EXdMuZdSrv+L+2fO0vOQGBokIo9GRGIeqO7rUWSzas8Xe
lC+UQH9uK/c878TZbqT219PDT70v9rXXEK4ThvfUgIS+FL7ZC9tUoPASM0rbZj6u6os2ISdya2CW
xvuK/nEhuIfg14PKc4KpJTtkZls/ux/FnNGF+60WPDL4Y3ClYnbzPcjIdcXuHby1UNGDZl6sDNJm
2MJ/6UU4hH5aTeprc5U3/Bs555jLojEeFMOSqM3kriTKd+ygIw4fOUbjFue/vqsSu8yA4Wswh/Pb
ot9nDahTjGhyPnW4XMooMXOd6m4F/ll92hyXq2csgyjeYNkmdrNJgFuc8KdGpQ9mAVjhdu/It5As
7y34VoZRDd9aKDRrye8B0cqzSgMkNVHoUBwyDAEc0+/dTHwnPyBqnDf3HJoi5EYVThsN8rjcpgCT
1CXoelg3Ma3vl7TV4m88bmloP8nQfWOBJ0TqHQzhgs+ueGvJvCy+Eue74LOnuEv1qH0SaQX5ywMs
rKKmxElPe8ySXTr6nz2QfF3KII8z1CRl/dQeKIHm+tgj18xlYmKR/Shr0sJ3Yh2XcFVNuUWIlArt
DwRLgaBbovAdnRxNHv68NG8hpfhN25fGLo4EqtgqzQYb8akxESkFvhQERZ8pqwEX8yqEIJSft6yb
dr5bb4pAc15Fj4IWUKls/ryFlUX4U/ZOV/2Fmflz+26cxl1D5TuOCFBrrzcK0+GBu2CSVXFVioxT
gGtn1ARyM2aUkm0R4UBuxRAxO8zr4D3wrBCSaRplHK6+iBE8CT2TTfE1qvhWcVV4poHlcn9iF8jA
C4xD0ZyvUPGYr/zEEtYWyHpvl1/ztR/2RLmNKkUgyraawM/UWZ4WE67LcMYuCWD0LbfUMxfFoYpz
kEMoDry/FvF0s9VrZzZWhfsUuYmfsqNKNdpSc2qjYvnQpAYXomxqjRiHLwl5fEjJO8nlkT8onSv/
Jdm6NgGVTyhI++/nI1ktOgPVm+IQRFmGgsly7m7Zs3ncy0NH4+RdX7+5wmWzwBlOhSKrqUl9lnLR
WMAtBBRyuJluf8J8qr+Hj6/YwRqQlP9kx9gt5o8o33kUz5FD81xeF6WsbkpkbYqkDYm0XcsOs8f8
5V7lpjM3hRM9rTOJyzu5o5rEuahZiBQ6Jm3ziGpilNMu+LqqObyB/P5N5ydrrLb2mZJUrdJqXsak
nAqHoQGY2JNOkFybWOU1pQfsDRrPj7/TQgtO5UsLTIggLHMV/Z3x7Bbp2q6wJKJAbJtV+/M9WRel
vxhx9hMrrHUHpgUUF/IThnXTYlAkVklh7oqY04BAGMcMGOIRHBdN4QJpdkpnirmDVuM7CyH2UChM
WZUdNkc5HTU5ox7NNKN9cjFDsGaaRC8Y0OI6MCKFZBrumpvee36t8wgqtJcEYgkM1+KJXAtnkMbG
S/QgpUjwYlgcWwTkXhQkIqqGzV9IyKK3G5lhJfhztVxpiQb5pB3sxypw0dOqOFAP8627llG//a9b
nuTNWojhODhz8Br6gv6lDgWcIz+ptqWXoIPpMOJGy51aUfDsSowxQXqRVwwPCdv5t3wd+O9IXX+z
qALTGfI4+X3cPrPIQ1OMqsU1cTHERbvkHveLSZkb5CiMxgT4qP6SI8xh0GobZEcotyIgiYfbFNSd
iWMdwmJ1tYnzIAUrn8tf5+Mh/d/V4kagLFep8DpyuS1UtwXzeHtqYrrYMBY/9oR/xUoX5UorVh/y
R6jNMYha+2eKPrvdQo3zUaES78Ghn5IxXWVi4oC1XMwhEWErJ2yWTPV7WHhKKdRTj99xu/zH8t2L
Mkh5lpFi8c/qdBqa/3+ZijUSQ7jumfDUQBbuzjjn7KDuvnB2OuDQxEDZFTPyfdMXcaLQwVQ75dHO
2Y1K396wrvJfXjGNmNRg9W403sxJKBHeQFFBbR+WQOOJBxCC1TH67naRFLvAYBcQzI+uFxQDypbg
r8QCVO6IDuZL+nj5kZEXSTkRnYeEvFegyyFmOWIF68yUuegJq+OeXgxP7wdUO34gZU8/pnGcT0Lc
gp4dxfokVnvtAwaimkxoMcGMFEXDh4x5fx6fc9X1+GokM8KQS2BVW6mfnCjXU7jWZzLN3LCjeZcd
DN/NDrac1H7wmguTlblTaogBbCq/5l7s7v3RMv12MDewJRAeH0qWDklDtmlP/2DdEZocPRsgqajG
BWYYF39Gry90jEw8dud9gn+lfrl+C2nRVfP+xteQXj/jJuOS/YKhMQRVTCBOJOqpDyrF8ofDpvGe
vgvPDwhsYPaw+VhFo8oJbke45ahto9sH9OVJpBRLhn8TGRu3J64Y5PjogcUzJw+ixmScSng1fv5r
omCb9jz2mEvgPd/8/zqlUn1AxEc6qtbVh0n5y/TMrwqDRYNPlkTMRR672nXTZIfJusl7Nm8DY9Mw
DLkirr2GcTOVSUFEv59lSyRqLOkiqWxL5toN+ssaxAGdimwVh1Dyh3YPyUr0VgcXqzL0c5BAOsaA
elkr62ADUsz+5S6NuR+MurlDqw7d6y2emgWieJuIVeS+s7rz6zzTFzvZBxY9+LLSHffK1xwavuDi
Y865CdUEWqolHSjkOiBy0B6dSJzLL8VZky9w8DbruWvoaSEGalI0ZFCukw4htoz0JFstXreKdO3m
Z41PB+U2+oGHu+8JeMcaLn795HT+E2e8hijMQYMXMzkmrt6w64P80vnzV8gPjzOYEFemV2NRnd9X
0cniufOI5vf5xHoxS6FaNBlg6wHLu+W8gkPrh7xhslQIgMr0UDuxZYFsCwZHscUsA8kV4TB4mkJN
q8M9uhB52kJvRA7Hqr3nNASdNXSrUCHR8FquB+NczrNE77NOQFOEfocW2K3tyOfCl16DWjVutmCI
jHMih5cjS5qGlk6EJ5CB6jiGo5SMh8Z0Jbq4glCABW7wS9iPCNWbsGJaCfcCHbFfi3eZGScTD9xO
zwf7zRi9vWbunueMCcz279nsxRM6tH6fbxo07vzwCdyCuWsoQC1qCtYoKguEAP8+rPQxg3EF6Che
JEXXsWScHzDiETR01+2kGDBv6lGcwDoYKkrIj27mJjTl7itVtPYL0q0GWuZwDYcDWn1VTlKCSI+r
3KM8QIxYTAyxFybOkd+XVJIfbYubWdkKj4WCGvohD4AaeDpC4KA3pbscHi4m9AybKMROgz6wUc18
Lxy4yq57fRjCC4Ozu/OxA1fbFB7x5AFKsR0Bb2petlgAEVckY7Q5XNgTWxJEQnei0IqW2XPq0La+
kLKcEYnZZgIvIavtpB5IW3fgxCUgxBYCPQw7ZNtfveTmf+HcyOk7Q8XQOiL5o8+bm7PbpkEdVUNu
yscuirvM748r6A/WuVZvZxPHID9vXvtJ5nxmMx+iln4n017kAbmIr/M5iuuRpbwgu6jwZUD3QsEN
VB9bx8gTphN7/CBZZYGv2SN3/KHEfVHwDToXm4C4NLJEYFN0h1RyDAMVSBgC7n3P8LeGsTq3jT9h
4joTOpxwMSyKTOtXdiReOxoFPfHzn9QOpL74nsYyBLEKjM8HAqcCLOhwwO4r1iT65o/q6KBRnfQN
4+upP9rVVX7jULuif/q4zzNByTMjPrDLHpTdqjZhSAlBklAE2swNissRxJwiGVzFDz/NpI56ooDg
iz6lA8ShwXTfVJlvINgjU1RSIx5F6K5Bf6ZeeCbFa0gZ3zU4UTOfewxR7McrtG2RaYBVaCoGctH0
aa93feHzlYLwQ1c9fzuCAAyk7GVswumCV4DUC7qO4FQMtYK82E7w0sozvK2Q4UcCt0WA9eu+UyS+
gLseU2++vBMZpx+T1dVElh/btdSU/0w9pC0b/DIFnFKKTB70AHEXUWrAV9Jjuf1VVo2nttB13TXa
Ufcajo6nvPvGSLou3kpfkCZxUxm+pvoxLH/A2U8DxEZ3fz4FiUAxDdPYQZufV6AM0iMGS+JA32pB
RZO3MoKsHy06poY+hIwm+pMEWqGscz/WXdBYb08SQZ5jn0kIYcVZsXtbvbm9qj9iol/kYzTAF1zU
mYYnL/Ggj1dUxm2bJ7M8bfpxkqW2B+E4xJTqbdYNMoNoOKTE7uszvpEK0gEH69wk6sW5tGLZcjMi
bztXdVNFk1VOGQhvh9/KXiA6+oG5Eap4/BAGCn4oR+l4k1HA7i62igYLQioGpJO0PIdGY/c42JVD
njiaOMrUST1QUQhzgmrP1j/fFLrGFh0XHOQS+snpXiHEFnvJOv9iNna67KT+jNFUiX749e0AEAH+
adF78q+iihKkp0pinz4ksZ16qGdXhVi/CiloyxP59UvR2WNmfDrQCun9rEyyiFhWIBXIcdntQ0ev
gKKukLoMsdtbf+3OVKCwPOZIL2m2bPFj7eW9c3yvCk9PrwhjeP9vmh6TyEOnqxH2ooPK44drj/Nq
NXOydZ26wLgqM8tr3OuudlzIOSBSDsECsKtfbfQ1Xn58nrIeZ6LXce3ZMiIbBMlLCBuEz/iWQ4r/
97iolcwa9Iv/lMD5AY7JgheYEqFZitjdok+E+0Hz3ou8RfDXK6VW6Ra68vbO/+TfefyOaXnFIHZ/
/6tBdz6lhGoN6FYtDsI7JbRn4E+HQlgegeTKGP0xn2Hm/hHRt6yd4MLtXpRh/3ND6r+7xCmX5wDR
TdQZqWJT5TXSEyNGBrCuOJPK4By0gXjHiaHb9dy5+tts63dzspcKA+aWf2YMdjtYQvNK3eVeRx8l
s9ssS5mLt9taf7Nl9/Arlsy8M3Aha2afps0GbhD3x/Tyf8ltIe39Kfb8W+x2FvkUTrLPHmcgQlIt
LGGFLV2+HdZM9SVkkoL1eJ9DGKVzVBss54z0Kh7gCA/UZxO7v22fcD9pCfUOaapns0FOuvaQ1w7X
tjDlQhM6EbDexr6EBF2/ubbDa5TNuUKSgDwTlAgEy1yAklnYcZO7yl6hWkgNzO0l/pTR/kcjhwhN
kqHwbqVejTp+wNjEI+8C3/et4CsNdFltIlzBTd8mTP033PPhwgEA7fRCJIFNIYCzjoj/BpTMmRlj
N2xpaTMCPYpEnbcAQzdfN4KtxGn0vBYhp8Eg759HDdV/sxA/tWSrgRptOkR4Zy1RTJav5V0LqvRB
OfI4rZpxL70eDncbDxz+VcOBQeTEBgLzZ62weZxQ2k/lJ+NunxEQ3KC/aP60RCTB9dtZNkHnVmiw
EkviYl7pGKmemWraRgKWQeZs0/0+Ec4OfuvRKhKDfEA9mxLQR//9/w5LluFOvDvVF/HGNSPdB/Cc
ytG0xxXw5R+6HBz9WndDSnaF4p4yTMCm8Tu/enc0a8xzbAh+e0wPeLX9heDjbW58DBGzunrBCxDM
wWSr2jl4LCCyW75fwxj/bwjF3MK7e5FBzH36LXMU+4d/YV+pWplnDhDr+4CjrLHUKF1NzOGgzTvs
7zT+vWiQUZYi2fp2EBML6NRc4QteHqs7tUVy+4HBoVhknIIWuG5QZdHFowIxjGRM/1BA4s4/tnlK
W3ZXFG3Opy7uptZomJ4bnDVq5VTXh0O9EtdjGJWGc6y7LURnGBfROrJmMXGHt0j31juivPJlKp8R
y+W4k0CNL/T9R7/iUhK24YGmm2tmu4kv6udUDotqOSa1Gg5XLRdiBrC+faX7uT6QRAO2RxTUruLS
RzHwk+e/AMhywolcDMTRaLAyWbChBWdYGrFMtLWheToRiMmS5jkALW49NyZ/7stHRWS3L64/ERwE
9WO8ZmhiPYdabEOUmYDVV7cTMZ/O+GWy0DM+9Z02NCvv7BtyhpMuivmrmI41w7C5zgFOOLHQ5tG1
D7U8dYLG3dQnXHMB/yo9PxEwikqnVEFoDb5kkZBkJVMSDkEh6iek/5R+J8fuOSbFXWK5qFHPltHo
pAJdQKTwMJgMPIREhCp6kvBUW+OVGWudr/CXaajg0Dgqw0CJ77m9lS/2izV32DMv8RJEW9d+qfER
5mQFJFn0PBSIhZszPDPXE+4J+9Y47H31B0nxoowxO/NTKjbe5ft8JzvWXpXFcFmUQd4vLMmmEVWX
U2eH/EpI7RKj8DDZaTzgvGjiKXgj/ZvuChSr3Zn2rrPjpiM07pt/njfQwIrnfxaUV4DLRp1TaUY3
kawMRKZ3rSi5XOhPa5jflmFjGSVHGp1bIS+eKB8KwURBTQzmQxoy7QNFGlzA/VTmvULtSTbI9yvV
tzaRZO+RYmDl/xbSAOsIZj+xPyfDInorinIeH41kMUFicg8RpAqoKn8LUDRAyIzlCU/KRedt4StB
luYFQSeBqMh0URozalBEGT4KEnT5WaSyUZ+OIeaT31qs8+VRrL2yOJSwWdS4WN7qLDZcJfwNDn19
Z3gNUl7sbadca94f47WqKbVkyOdEOADu0cf9aivG/nv/vYbMfk6rumROoCHXRnJ0hu9HxVVd5/fZ
FtLyh3+K+9kisQdEM3wCqSKx5PeVbLobozDp0whrnCyyVICw1Jr1z9gU+QeUAVPb+coAru936Xcn
fbLMh13qdZvuUT3QwPIgSpKd72N0Cn+nAFURxeXadGEDbI+ThZLabbYo+D44b6A8XxsHpHquh1BY
bA9jttjNXwcSOi0FdC/yuv+1T6+PqbMW27r0AdD48vL6q6H015Y5N5D2mfgQobgaRDvq6gFVAHwR
ug5xXhOdVNfKk796WkHYYoWKZVMCFDg+lCrGfpGWtBJRPuN9634z0AB7ZUpY2CRTKcRRmTZG4BXg
CTbTbWC5YVI+ruzl8Fp7eHpcWjQboiVvCVTTHw2yPr2I0RllrVB7V+hbE38vM2ehPPgZkwKdKFJr
0uyrgWdbxBwG5tBUngl2xdgifDCoyP/pnNwmqLZkFEm23TIkZ00T7bjhwRZfZHjmTCAQnm/RKTcZ
J3KralqcBNrXZ43d0EfqcXfPCugaKQlHwvct5+MEqSO7YojSz5nI6SG6OcxVmgvB5/0p60S5W3Kh
Ro5a/8xnD1nyaxBLmiyoZ15MSOuXT7otCjZgLfORux5NomnQar06FcdKWVedPex3pJyVU7jKkiZK
L0D20pR5R/Bxurkq9KaK2zfDzNUGrRJflSJKGc0t8dPFTZLa5J52q1LAsG4RGwcylRLF/i/F8C68
Tgsqjm/h0ODD3lbsmjazkA1cV/lUetOFbneff/WvO3acI002McCfAfDIJHIgnylCwWLh1GPLz3l0
b/iPzBhvzYBldW36d+q3N8w4q2ja+Ldo6ZcWRackrYQ7skY4FdvBW1x9DkmCjTJkYTooQPFIIF35
lF4BkrSE6Fc4lVSMnvxiXHINdQeKAQYC6vNhD06sqiZi705Io9wfHXceT66zGLbytR6OXyqH0kU3
LzTCYpAdx0ObiqoGxSqAVXRLqFiZjp+R0Et/ZqyL7vMNdNrrnhS4X5T5AnDnF5Dtc8GmdJHUjere
MBp8ZIJj5PhSwRRnVCeWhfyK8LHTXBioHwkGI6W1o9bdKjr6uvjfT5lklMwj3DDAcdkfzOnq9B0a
ceMJFAskZetGQZVxngJyYXR3VirYBajpY5aVIsdRCk7fhn1tvP/TcIPV9qjxYI74nbju1irl0j9g
I/X6L+8rQ0sqUkjHHM9ZuDsEv3fcvnFFoLTfreqd/sLWdwezb4wR+zlLVW3AXajwXhIdLNdc6CD7
2ULDZ1v5d3gW94Rl2C6V6FQZFne7zvNoq432q/dID6WjOFmuAwUqshA9SwjMhjayPdPZyKM0UQhg
8RcQR9atQE/snnP5/XMko74WlAR4zncawh/eP3jPTN5mvYthGbWs6IoWyaFyvfY+lEOcXDjp/0yM
r/gMLBqdHyH99G3/n4nZLze32jdgoy+aa0hCnFFJFsGeRqMwP7U30CPagiLDUefs3zZpxLBIUNyu
0f1Bd08K/Z6rd/SYk51ESntSEefbsKodlmTElDbDuy2ySlzWUj+kMsK9JgreSohQmy9rXQoGbY5d
42QIZCkcVhPXbu9n4I6wX1ljzj2spSnbXOnKJB7lYAvCfUeFXkkqYd9GX9LWQDqFZ0MBsCWc/Oza
hUHm7884Jwxe+P97TpGtxAg/fvoNYNwsSM1p4+wr2YdlFfMbMm7LlmUmFlsN+TQzPXTkDt1TkEYi
TLl+Wj+uMNY9cylKQ6LEQATcdztdxXTRxIagv8o2gmo3iy8DuT30JuESo1JPkzxtZwIEMD/MVvOY
c325Xq/ZV59/tGAyUsKYuaaQTYybc71hop9aC3k2e4B1Rr+GkCfTLt+bc14mykDzyt+APcoIAKyq
l2noRwhGkzR+VowvwAsrkaRW+Vdk29Ss5+RsXq+wr/iVG1eVwDeNZeHel3QpOlwlrX6r2jYKeevL
1rsBFuNIhHCQAxSaCJScByOIwiXnlLvcX50stZgP77mtugrAMyL3CNTEMxWzp/ts27UGqVMIMUIP
/wRh0l/6KeCqD0jHEd29rxOzsmXQsaWGk/XFCYhhX2bGteho+WbRAG0CyrOlFskeMciIIZslBenA
w6J9H1LJSbGZh+I7Wp6Sj9yWMmESAGN/s1RhH2F9g8Uu3F035BhB70fOqiVmPJIHpPq5Bmo71k4d
qVILzzO90qWCpYfF/0MrsgiN1CuZGWeYOI/RFtDgRscK5aCdeqigsP2doDtoRaWUcxiUcKFjl9PL
oQGabvyPJF5znQibSh6zon5FFomtdODSyhrm0lVBkAuPM/uzSXjU+2g8UXndE4m8NIxnN1aS5yZ7
cmdmpccoXaMGJHjX5dExtI9h+f45FNVL64Sn/y0VmQgF4fZRUyI5OvMW5NKCEeVH6a8IHVmoRd40
eu48EyjBjK9CVHszRC1DY0Kd7doqiw2ZzlgAkGExcAKOWVjicMDD+LPo1YNWqkaAP+Ydbj7RQ0Cd
o99ESxjmBWJYKovNElzPenkWDaivdGkz9Z8k6WRMGmJocA3PV7UQBWZoNwyaM+M/fDEs4rquBQlY
Liom95VX07FUg/qE9erZNBpGMB0zyYlTs/MtJ9f2omPvf7B4Krz6MVJC7Aq4GCOH5+FY0aulH359
UszTk9L5zsjd/vifNsYbkpr19hPmkpdKduAiBHcxnYVT2IEjRHHWJH3SBgll5m/q3sHSplH1sl3U
MuKdmBUw14oLfa5frNBr4h5ZJYliJU44Oshwe+u4z+3TSVmjRE58l7ewLjFua14OYoCQHcldpKuG
zm6xa/l8cHyBVq4UJxY8Ih1QZBI8u7lDK29WJ7jK+zADJSrMAJrWKX8/dJR7GBbG3ZHqfT26SXXV
9ehv3NtJYLywriyYKfHaN6kg6ynldDcZR19Vyg2bxi8sEfsYGbgGIz47jmcWT82odSUSRG7HLWKq
bd7lmlobM6dP3ppZIvSfrCgcT2V8VkkJrhj6Xa7cXwy8mtZmY1/8PIpCof86iDm+2aOdgWsW86Mu
u8lLm3U02kbwoa6+rnjRQ0BVFJh+dJ4R9jJTr/prZ7zsDlXeSNfvB763N05+CseHZnAnNevHl+18
wZyNXAfK6GxNLjU3KYkAadWUglpKmzNy2QhS5m74sG/4mgtxakV/ZemdqWy35I/kpNP5M52Lao5u
aL11As8xjfaQEggxKheHmEPPkeTwz88QYNJQduTa6u1GZP1nA++GbAvzKsT8IeMmfJhZ5cAVDfSq
P5tkmpksKrvthrl5qcK86epKqRkA4+HPMcvETt/F39fplYarQZkBuviLd6KAzCd3WVh4h/qJGHPN
4f2pLfKL9EhzhvtJygm3dMXDgu8GwPN5pek7W1B4CRvqeHOUwk8PuqMTdckmtwKPXHlap7R9Ym6f
geD+M0nJz8rccfN++np7sEc8QqKxBxThd1c1MFIZIiXguUmpp6/YdXdKSlsigNws5JBHnHnGHqko
4m5su/s5uFdy76WFT6/D+L90Zu5lytwMtH2nei5DifJfX3/JEG8Nunk4g+tIhyBdFbdo2rHK95mA
do5OT+b72TR3jj/dilFZFKiHkOWssb5JtSUhlb+KixuKrTGslDpWd1phIPQHpGRlKKkymUHWhD2M
kION+t8gmDRji+JoOV2zLB7/Wv23p6RJcnxetqFXFvMvzz6XO9E4/PKTorVtDnPVZUeggurU3ysn
+27egGSE5ZSm3tsqIVzXNN4GyK26TvL+zUbazJpitv//pTnBNTmZAUSMudkj3v8/4auxhnEOCfJ/
aVU7ekvf04anAxilfhTL3Aeq6nVpgFtvA25i5ZF3r+hGvOmMEFWlhkYKFXJqVfj/MChqDTmX70Qv
5ZyDiaO1D+SubiXNAFYgV99uGjeXc4eeYjVwStMzNNY+qSlCt2R8n8QzCKrpnN2afWHavUlg+AzF
lVnTFk4OaPCMGS5Q08LGwSxKPwwyviuy274tOYlU1pIE5T28DHlkKGh3R2FER9i1UihKNfSvoLjq
+T1/xp/DJlP3Bt0PxhW1tlUagMfcVrwq205zMIyQs8eFj/TheAmVj3YMQNdRSICRN84bY9/fBknr
2mTeW9DDKOGmYy8+0ZS0HYsSNwNdzRUSyO/HkhBrHKSxSUpWVdOfRtd6AhHvZP6eSai3Y0ren6JO
kr19v8EkrKHEW9yuSVtExwOXsFbicvI1VdveGsrlIcpIpxEf95HQploKFOeScLNZlSpmW1DHsi4t
i6izoiiREh/JAPBTIP49SWlLdeK7BaU7NDOt3/708bmjclN6oLpZZHu0nWqoQsUkyfZ4DY/Y13c/
lb6zy+y9kBh83/70irBz8feYo8BIgBQ9m6eoatYhD56gjMl23cVKhHfU9zbxuV+V3BYafnNyF5fU
U/C+BXP96+LW4nvM9IHnte/gPQndaHMNhhO9IU1gZFCVByA9efqho71EsEctFIdSEOykl5ut6BJt
Ya9kcsrWZnleG12wCW9V+fVSl8xhDwPn9aI/LRbDjwXiARCC+Udm+06tDA02OWJRentFtjRvbmcS
hOgkJGHqu/xqP8D1dfbF/TSV/Fr0sgC633ux9iv8k7TlLJ0ryUOST95GxbqKaG0UUm9F8HLv1G1y
aEen3WuYidJ1kNHpiqUWBhO3tDTipupUZxh4ap8UAuH2wNwP84vrL84PyiugTLaxZaTtLxOnl2r3
0V6/rfzw8kqfd3slthDDs7c+SYcSHsoFHFYUIZ4X0FobPasA9x/j3zofTWjLWh9XHQeiMWnEWuPx
ihUNHVjjWE0y2VHJvb1U2mUEoCMvL/LxS6+4yve89SQaGLhy4YptXdAHs5dz7Zmy5H5CQAqYyzNm
iQXF/CrxwzRVUYvVjhg/dy0nJ4ZcSXHgPuDXQua26B+qrFvOTQlUKsvgZv2XF4vxCekfiEh+e+KF
IhEEBWqf38CP6pqeE7aiJNUnB3RBFxOYdwT+Hh6G/vq37eFZd0fRZ3AMQZfh1mzX5xI2uQSXsnsv
pIisc32IuQFyfyV5ERCQxS2Qd1r+WT9yVLcWgIu2wPrRSUpM6KZ+CJ9HRwXcOzZPvZjB5EfSfP4y
jdvHGm4Ez9kTWAke7eC2NYbUcKZ4ma8mYdE3gM331jYLJej8sZnjPAlWMzQloAWcfLp7O5KndQd4
tX0PIANKLJ212zTXKwnFB3lJG1q5tp3Uyq3QkvFlPMKxWSBxqkypHYaANyAKFGfsn9vTw5XQ4wYg
jT/p5ndaI20KcaYaAniy88te/sEs6zndGUVOg88xP8211qQECQOlJcOaBYqm+41N3t3bDPkX1fam
xhtSLaCGs5UrCjIU8rQse8soDc4Rv2YfDmtMJhCc3+s5VHP656S+5fNyYOWXHBeVqATXaa8o/St3
az+xppameeym3xPBvKG0l0cA+yKNFcT51JHls94kJRviKW+2Y/VN0zdmWqZF3x7irsVs0xz3L93k
uBJjFpiL5Qk1kgvmZTHCLZVSMZymWQToaUOnLenfjOm8PLwKr7oHKB1tp0ggfe3nGwLmm/Vvp4fW
g4GBwPOJ0gXWqh7G/sLus7sWQBF/qX9xkg6X7ME3E2kU32EjZcTahhDUnCYZLB2TN4BSccogEW+J
U4L5MMjm+Cg1Nge1xeOmZpKglofQI8SWYJRG/46Q3+sDyOJ4boytjnJ4YnP7bueJHhj1qn/Be/Oh
DGGso/ag3xNGIG3cXw8sgnQ/fUziIQ0DXhS8r9xnwz10jdl7s6MmQtyEvsn9H8bU4QAj40u/Poe9
++CUNdISNCsk3Si0CAEe3wCyepz572adAPG6ZgNTfdOOu9dmmijTOAxoNt/U+nufk/Dj+C+M+jyB
hYS7GQDDyO3aVdVquaGuizLUrv+MssX0EjglcT2vvd4BHgtAoE2sLWbozgWingyIw5E2qMFAVnqa
eZCdo7QUWWhSiaazWr7Im/WZKPInt4ef0YAJBrDVQQB66rpl9FGI6he9QXC2snqi++On6agc+ksO
MQ0LEpi6DBD4SrxQmdp6/KtWUystuzrEXY86uC9qWeEvkQBrmcm1Qi975qhjYGDS4A8D1ZdG0O2s
roWXWL7LpBlcNcyU2F4pfFT37JOc/+URkVIa5TXA8OiVrAUiEJpYYaCpOquNk7sVWdkHA9i4T0F6
zR9DqKX1TMvRX4imM2e+GrwcyUp2kJxPlFWnWL2a/DeNng03y8DXmltGjRNO4VNchP66NLcOMAqy
m8DD5OykeYhkKUd5oFdiWGKuZG1SD5jWNvNGNxiccaWM8DPjKWRVWfA6BZC/nwyOc3ujXpqPySSw
7GlJlZvLaHA99tIVZeejKcIj8/n97kN43F8RBEVsIoFKQ5oisJHBsZg9L24wvKGCNJKsJs8PwOID
Uj6iWZgAaAgE/rq+oWR1dL3WUaLIcW8KGXmJS0RlSSUAlNWmrVSQ9DMt6l6lTMpyXMGNA+wsdoc/
k+lWrxd4qE3lIjoFZZqoDSDjau5XkePG/D7eceWJm4KtWa2qDWKaAIz6tD4qbAfSdZEfO/2XTqAM
lVTuDR+kIoko97IPcwFSnqOTsW2zEqSHOlWjfTdYTPLACBj+tKTEUcTrcyM/oLQjgXWam7iQ9rnL
hC/M9VUo3DNXYOgXJy/fTVhZE3mfwzY4M2MBPnET7DHU7yZF1jfs2YngmnpDHfVQxqOc39cLvzpf
KhlIq0V2Hxevwb7SI171r+gVKevIYedmIKsJCBsekKWzTsDofCxiBOq8Hwb0wzl5eKX99fvZTGQU
k4tv551WHabIFvUvAaVeXaZHboxyEYYha3N5oWqE9LB2vzmAgz3FA32CceeL3Zmenn43aWagcihu
QLf8QHKj0O0O9Dy+2KiSLtPYJEsPvsbsJWe1JRfDnqHQl1uvualgXegBF2lC7SRkQI64oZ7VnzjA
kUkO/qHRnmqN/rUfw2PQ8v97/xXrqGCqx2wkc6wr3H+kGF8a5ddgxDnZK69isa7YbGKC0Vv4Y1uU
Q4NJOUdk8dBEJnnS+huuCdseZ7cZIfpMY0TWqe5wFtVT5ZSnERwkKSbOh89d5ddu9MukDYquC3cT
5oIZDwuFBHjcTQjrT/tmBuAxvi9EikH9xKDs0seqH3tA7z2S53fVytgIi7CFCxXaKrvnq+pDJvQk
nA8wuCXMvS9sKZMPNjKtyKfKaEzsSxhdvzEGACVyEh2E7meC83/2KvyXnrqODwAMhu252NQVJUjW
/aCPUc4fTTRFLYhQ2KlZ1gVh6g16aFP3mbCOVDSSXdvlH72YqqtvmpxzACJrm4/BMSX1t6t0/HC4
yGtWYQ5X4tjdl0E3nzUvCF7f3CkGlca+5AbLVChJDv3jNdCWI3toWYY/+jdBzv1KRaZfdcSRF0nJ
2rGiDHz87E438lIgNGCm6P53KOD04MwQwAMGdDpC8jLF09qnwWFKNZlYx5DxGuqMEOdHquCorcLb
9IpJdTvhZ0xCd3Twz5yKFxTvGDbr27RGQEHYIO6jyfl0Igqq0BJeeb/RAWK8GRfvw+oSr6lenixL
OU58lTpq9bk1qkc+BFq/yMFLcY7GfWAblidN1mle6W95w2eaCtEaTT3MflpPYSZZiatfvTGSAbjN
6rxnetYuFp/9Z6pLIVJmsOWAhARpdmUz4gR0ubR1mesXBBEi2rMS3wztpDEfdMg4Kd6ikPhgghw7
BM8tC+BwQY3vrhTchiqZ3U2g6rNVC9QORG3Xoym3YVYIJ3h4okJe+CCbZUpX4xTmcB2DSQiG+YeQ
GedLjEmSmXOuEta7nTLtya+PUB2EW3iM71V1SxNi3WZW3r8BWhEWQzB6LOUZMuMBa+fB8xCk4eBD
X2ERumADk7p+KcTc6F35RnPlwal4XLUqEyjhXqEAPtUQMb0uLhTwXH349vhn9hJL8AraTCGggW5D
n9aM/dkQ1toXl7mzgKbVczEbCq6ruSW03ua4LywsVSreXKLBMa0AcrMngQtreYkmccYglG+Y9xNQ
3wZGerm6OGsq3psHiiYXGTzueptXSFZ8jR27jwEftiYKN8EnItZABSf+9uII3sgryxS5D20SbHDB
xiVjOT6bi37vp22I5AydA9bXk/BOlyuTtcfpW5gOx5rr0DiytBWz6YEy9wNx70EBnbbsJmO4cAx/
qmREipatt/SV84fuq6m51VbhgxOpUjTz5PhowYOoMd1Cyxomt6LJxU0LNWfo+vZZkoJg03rPSqAT
IWClkPn2V1VvtyPPcvjgeLQcdS/hOknWA3V2MVSsWCH8hCzal6MLMJysPG1ME6Y5YQ3s4/qxyxw1
3lvESJhqCujs2rudizf7gXnfbNBIn0QpwZ9HalSa3PS3fQhABTiOSmUec46YMN6TZbdGdW7r1m7t
pSZXzr8WqI9/uJMNyJvrVIgNyhzCCJzxW5j1E4jXddbS1neObGjBHPd4cM9pSzLO/q8sybB/R/G6
S+trB6PLVajmC4x4nNoS3PJ12Jo9qdrnxXb7uuE3QL6wNUfTCfhW4of6Iuk9zESFSpWQMzQ1F2I2
9fk4KmS2gkKadIMnco6D6oNf7d6qAfmmvtqNmKuAbF3L+owcR3ea9/oMGcZSsQObuLi5OHjbunvY
LpVtEoJn+EPvNbmvzwtVEDn2PmtNIoZyKfuHVc4q1UfH0AzOiQk9ArYtAdjejfOL+CJSmi7lcb67
Kj36Z2yXVWztXa6P6/s37tJSamuJcrW41qFXKlPaAf+ABNR1E8dwSZoIps4cONA9VT2UWtciZKwg
cwQBsvTXTLR8pdkxTvi7vlw7Wem9TR+0K5PoKir5LYvpJhW9+E8YSRY4ihEfPJjLh1rY5p2XQkTu
z7uH7+dLrifi2H1+wBQ6wzDKdOXW2P08HGLhqAIMgAcFRh8+jSZb8H9gYc+MBMIHmfaxny/GC3Uv
fuOGhzbepwIsjziFS6Aqx7qnY3wGSXg4asbSsApQe0DqYChqhBTk1ubE1u3d7ZErFh3akvOQynD9
ICu/c6Qq9biAxc6xpD7eXtVUWYtelQILTE4KqRfgRCUL5x0sKu4DQ2vxwUxKU1txATOsP7LWR+Ok
q5+nxVX1hQIBZyRpSKFH29tH8KOgvm5Qy+a5RCIYDbj/QEztaDqXGdouVNFtQbuCQ2tw2QT5AxkW
POY3w++ceemyr/DDjIXAEhNaRynkK7n8i1oH0XIQAhQBnfIzL3/xmMC3BQFaSh7vSSZ+eooGn/65
ks2rj0EY8Hi4KElHp4Ca3eTjdYpYhHUoGhaIWuYqeWHIdQZ8FQTZK0sVbMhEOViPbHhA7esoQoDT
1Ma5Hjrydt1AwhxAOKpCNa3upC2YNnTihHZo+P2GRMrjVEJp856wlU9Oifl2sOOJMSglTX2kX19b
ssCzdX+wEuma8B1AhJTnYpRdZuNqRUAm028ZoRXPovNtXHk51kHdRg8ph3nvzM7ZdFjIMKqcJTKX
TbQtdHQw0FsaWrbcnomgGYZ1KoNI16e+/2l3wEEch+/3ZvMrAeD+YtGgcjxBTKe5YLWDTYR7tf/M
kkM8GeoqN+ke5agaciAl5RTo8oalsoptyp8+XssdGBlD0s8ObvlSRQAOzZsUEeP4XoqqMFP5tRe9
j6Bt8u/wvNK4I3qw6cmJMxSYCPCiFFNYCPJaN3DZA9uG+V4rwRYWAwj5TajvxleFeTDKcuXUuxI+
GggeLZKamtz5HoVjBaVBtaofKHQVAW2dp5Y83E7bFYTHH4TnrIZPPggedttOxsOgkaRsY59KLm8C
gKYzUoRgxnx8Tj7gGnNzAM+3wEzKxnorEpjzQ7DMaMI8KlZaO30/17RmghrzT8OIYivngZPVmVIl
9f5K7HVSJ2eJqCyX1cmeQ+4xBef+AAa5PxIQY2AhwgiFSCwvM4kMZng+Dbg2Pe2qHDioSzI60y9I
FhoSLu386nIPxqqr45owPOeILIakRnqLg3zFAYbtllNqsT67ajqj/gCXc5rXCjDPxVh9wk16A+PM
t80bMETawmsaeP4YRXLgVrpY289inVGeHhJrZpSsTWooPuKqix098OpfZP27Rk68XjHfLCVlV1EY
pStQfjgteuovSvaWFRIYFM6g438kIBmm6f6fN/WJPbmCEzBc47H2IaSZrBsDRU4mLEem8HGiQFq8
jn+xv7qVJTa/Hg4QovknNeBQU+FyYJn/WJvNQ/Dgut0x/mLGxgUzTPiEzn/nDhha0IFc3A3VoPkS
Hd7jgLLuBxEhvEHhKNBn18dfqyNyP9/Qwu4G6NaLQkGog0DpCvgSxrOB+vd1ZJTRkLO41SuXCMuT
xfuuCFMaWI+ggYnwPjZA0HMmwO250HchXjvHoSOqN8xFG0iERnnzlEe8hGH+lzpSlDQO3kooXoJL
5s/L1DqSrRe6yXjvzOq9UonIVj5KwNV5AcAy4OTMb0BY9B0/LEfkse54IOUXZQ9EuSl0SyWE9AH6
6a53wnNgwKmjX0QTuJYKY5doOqPCa8LDxe5h4BsQHhS4Ndeabmg8bs2YmuJ7xrMsEHWmfo3du8WW
28ME4Cew+XOiRPVRyW7WbKuky10449O8qbnjNj39unBUtGv5SrzaA/jyxwcILOSkzcqWIf1agzU2
+Qfwjr4CuqW4CEwh2Wgo16yV/tByssOlpbBif8Q6rfNyueaGX9LynsV9mqmSQHRneG8w4lw4yX6W
3Y/q9e9YnfPznf6UmvZko6qQ5sitt9oURTQFTzVSxPE4gMQKykaYLxmtarBCGMpObGzRhpdrFMaA
YrKmfkdeCT98I7yhikDnvRZdsfRpaRdMxhiDlbnyaEcCH0jTDCrINP7Zx5NYAKZZUd/r+H6v5xKF
BjKcvSepFCibxCcpPbPPiVJmhPtxLL5qByeaYW6GbqZ21ZgovlqVOzLC0wyBSc+Kdx3htdkQbS5M
IQgXxa5tQQf2r+2tZsJK1/jsOduik5klnads5xZbVwOYzYsJxD06PRBxve9tZ3zF9GCgmEdZ3oN8
0jDzwFizs+fyPJMEgVR4VPt6qkonz1J+Cr+YieRXX0SSI+tAtaW5sgTlVoU444CCmZ7IrNKgxM4K
o6Dmf2VbxLEDcdK9RVqAQOzpecRoDBa8p7Qhknv5eEzf/zwMAfHrnNqybYeCrIW6/358Mey4lhhA
V5iiT4L7GpjostCA88WALl5Ghc4OCSb/ZVgkDJ93zNG/VkQGUlZkTfll0tnE9bcgNANy6U7MgQP1
ZZsWDt19l000AifFqwHf4DqRMZ7LmoEmUH4E0KdXmYHtz1Bzj3fLZPEBX+RN9h24lIDuNnJBVF2M
2Uk4jddKMAk7/0N4wZw8EH4EUsSvEoNhtzQhxv529piJtKK1zwBO2pI6PdwpI9V7nncBNq6I6cgP
SE5Tp64CKjb0pYI4T8kwlRJpQq/JTkeGQpSYEYkNfHuMFDTcQDZC560MFRrB+nZ48udbPxtQ/szt
l9bQ3aSiBpmx5vKccuMmMbb/s8FFx6f9xzYgab5D8Hb7WBE/t9FAgJULNC2UgqN3Tg0yU1J1nIK7
5C0Pbc+E0M/w55XoUiYSvlXgAFn8IHhkROxYQWl/Rk07ixVyGeXb+C5juNpM41wErCMj92ZyRLww
QGDQMqoue5o7Zb2usJYA0I6+sj1Q9yMAOe0D41r5P3y1TyoekeITpU3SmZlo6C1tPunxfQZUZGGL
96XrtwjN0SrVJBs9ZT1vbAblA3qRV7pNucjzlqjLwq5JzIoul1GwHz2/LPMSSz92ZP541VJSbB3T
qiP34TFCMiugMUpqy/Wj1qDTqTugQy5T2K6OaPxa0YI15MmNQkv+z25DA2F4o7LljOA7MEh4qVe8
tL0MKA2y9m9G8d+T9JQDL89JwLeIGdirZx7MW23QxyzIzu8iG1SWc5goJd0v50WyQZFbOZVuijpW
O8zoZK7G3IymjiVKi98oqHWezHdxz3LYhM4wy+s0BAQBaVwUHgIQvken6UDocxVxqqbNFOU651l2
JquRJ+qzXktXKJrrYnM4tsdeWNhk0QST+ObAly+NhtTt2nZXRFvbol5oY0Ph26eUVN+iQBQSsVeY
0XA95JeRzsC7xauNYBpO/X9Tapg4sb7KjslzaWTpY+HzJHwWWOBP+VlAAlF0ClU4NL/CdLEcljwN
A+YlTDiiwj6WhEPA3zPtLGvaFFxHA0tl7ptX3eTATzQwy0djpV1InjaDgL+K0CF6i9/Ywi75Lx1W
6mS8SDsmQvE3HKxIkV3nuDb/hRRaVNl3U/Uunodb3ebug0cxV0ZTcGVRkwq/Dd2XXl9UWvLqsA7E
BxqsVJgOMAzrt9Y4G/i+n3WECHmaSg2jOYe+zlUr5EBWEqJHLqNDZIv4eEUI2O2VgF4FIzrywupi
j+6KXpeyLoUGa1w3EujbP2JX3s68YFXtO4Z49n7QNzUPkS1b+w1vmo+CtydR4UfxQF8Wbme13KqL
9UHl+1E6/zB/rhXeqwkO3VG+m9sCGWA/+lFGdC/BrOUetetOcaiAFHuzA65nkt78R52zWo+L9QUn
5Qwc0vf6oX2Ch8ZIT9jZxSi4NkT4TL1RnoXtpUiQQta0Jw1tPDbRNbpupiWi5rSTFOa4LLZCise2
oJmegCEOPzGsVJRFWl30A7jkGGNVg9m1a2zldW3lh92tRiRT/LH7pc/y0dOkxnJCtU63WyAJXx3a
mtVNBTlVfG1XXiLAg9HOAyLWD+q3eBDV1mipr36tWtq0ZHOfLqNXk9dodb43sL3wmrEZIBYdatk7
ZDpMMy7fty4wWYEZR4iyfabb2AhBoMYT7cUnAKveOvTzdG9/JggzorM0VTGFTueEW4x+T6bMXHYa
JdOsOwWVCnIV3WEoDkfNoEzJpRNlLjkYW1NGPxbdeacl0ekWeo52hpJkbwC3lNsu0IPS6feXUJje
HdGXLpRrRIF0SfzTf+4Y6sNGb/IfzXGaGfQVWtfXuVhw/44k7EpMLT2G8IbiiNg6XwOhhJSj/TBM
9XEQGMyB+T5OL4cOvZIkXojgTHa8JE4yps5OviNDpNd7jjhyI8Kao9tWTmF2KTDj1FYGZVLTm5E9
nXdbT+gocqt4a8MEzyqZpL4cf2AnIvpU/JUOovB+uwNwAHGIUzubyWFiXfpWjomfeqqLXvmwuyEO
IdwjvwL+Quk2bc1niimaHPjgkDM+S4ho4++Ol3HvPTQxRYGymhhr0YZbY6Gbnw0kE1piAIIKbm8M
C6L5vN7Kys8CCTfqcf6vx0oFw1MKU1fJVMUskbt97EhFYG8uy9oW27+utc0/P9b08jlVuw3VQCG/
sE2p+n/5f/Ga9wbZjou+xY/HlQYQkqk4UU2I+9kAde+BH5PUuzXYiXYDl3VAOUSFHGds363M+LcC
Px2xH6Xdh6yKpgC2UNcYNXSKAdqzdCG5AxPjITyeN3taozwgO+hvtv2TqHEQ5F5LtAEy6T0n5U5R
Nf7CuU+FplPg2pgJoSWUB+7qG0ifugaQTx2uIfl8P8RJ/2dVkFNVCnj6j7HzLNxwrC2DNe6sA9zV
6XCF6DPWY6z8c04IaZEZXGGJZatjf8Lnd9fIB1PHru1J5l+yO3NYrpfliNCTdlehzAMhKIaI3tuH
GftWMbW0OMObGLl0bSCGOgi9z0ejHJ8AbgwM41qw9pXCQGn76ncefEeZBRZHTuBDw0C4zBVTxaXN
NMc5W1xy0TTr6HwVM512Zb3YDFL460E0Vzbq/XMXtwNldxrsWmqeVTcjauc91KBTdRoZoOkWTnmu
+yUWtnbUfvlypY0ZVixGBiwJueu3ppq6ccCBiq9PswbhqOFrytHz3fdamRbFk0fLSTaRfainyvi1
4Af0tKLCYls28XYm8KPrE+BFiENTQIYMZ6hlVjrdi+8af3pFVAEFQnlPTYLQMapbIdnfphUNf21N
UgkeMCwzvPZf1hI9q3E4B57uPdYc70DMeP5TLFFz94kDiwktpEyLik6DJUhXCXTIxDcydqF/r+DU
al9YAD5UlZxlR9dG0aGmk+DxOCBjjxFZVIriJQuyVIGBGpfTGyUlCA8eEYwyw3XgkEPe0UA6ashI
CM1jMFVky+3FNPo5nBb0g1p6FVJ+IkIINJrdNKwx1NF1WHcIJBHhdsuPHWka5Tzw9fvbnTK6ZprG
hW1PtYMZEuDpUyjnGAs0+78BpEvkqRJGIfuswIJvNR8btubogJ7NN6G1zj3K30W+N7tvPMgzmT/V
XgJWrvpnLsPganLIc73ImJOwVDGUSYsRjiPBH/6MYmq8F6dGflbKWhBWwUvbhAPZhsILvB2UiFxc
9GVlP168EH4q6NqSfBx3zIuYvyDX6v6QsxzJVwovHYPdMd5tTRxlF4a+OzrW+37K4Bl7Vd4DGC/O
FdEfgh0B7YnLwAUZFHXel9y4e8QsNpSY/aE+R1ryinfpH/lr0O2k0L3w/RNGkP6ujjZWRajrMVB0
KJCOj8kTkYv9KNFVFnJ56A/o5YlfJgbaVWxldRIt3U7142M4g9qkxPNak7ntm/j2vyME88RSsMmQ
XC0u9aLg2F+ZTQq8Hg6IL3slT+hpDOM4601Im5VDGPD1Cko+Xq4wERneXj475oXKDmaqj63zNeqY
lAcXC72zBSMj1hNewrkSprtM1vOI3YUVAek5d1S6Uyb2is51zktqXg7be78sNg21n+lUXBuxE3Rx
zqCOVdu/sRaywNMkCjOeZ2FDQ4Z2FNcYqao0zGRg1UBWrDnC+5Xusmnhp6UMmhyaZVP0iT/LsHeH
UoTBXQajTfCWe1Q3Mk3yTqitrctMzsy9ygSMksleJTnyNrKmlL/gTpZo+LSBUwqlrI86cYtGOIK7
LpEVsLrxBYW1/jbhtmag+9KXFu/GrE7S/j2XKdsjM92Gl4NIX3g2MJU3uZD2T561v+OaEzdgpLP2
SnVqls+PELPwEdEoqK8iWBI5os9EcQuu++8CPOsWkm3sjygSZ6ZbN+kydNnBF18sY4M9Xyxm5jcU
3Yb7xC4i/BT5eJsY8SOJ2WQcKr25h2ie9n6gEryj7Wgx7e8NBONhkIF/nwGZPrktS6F9kNb1vyQm
zMDNPd9vXCpk1EqVHH/fssXo9o4YVvqECSFmHRuYOVQpRG2zyaEfXFC1GC5yFx0yEr99RpNhkdnO
OC0H4+pYTZeWuRBT2HPngn0zdM9kBxuIlAE00xakH+RWzp9qRUtVua0mL+gnMHxgn/2WRE5Pc4GV
A2IDOzzikdiUR4DMolxejc/Oj+LBuhk95A7QZ/aybqoI/2MhdkkThzTgpkPtz+hkZfUmALJTLnEF
vU6nUTyU8vABClZ8aXVoA3fwnOKvEZ/mgzG4McRds8R8Z7sKHXqOr7q9kUh1EB9kNqoxyLmucuKN
BFFLXw7NfsAZvHV1QbgJKySrE6Hnw/NDL5xD5g6TEUEOIsudjTV3lYgUnp8kPRNhQyyTzE96Gkn6
W7chgY20q3oK08dfvRBJzxUf2pFQ1sf8kxo86Kk0hHV7ZYznbh4Tgf7bGXZ0c3x6RWOMExvpYAED
i7FWuwh+SNHNxHoJK4/p+5oBhwQNTjGbmSY5j0EZz9Ou0KFOs8WFMfh08/3E71rs70owhzwKPRWX
mH3rkoSnIay/RtgC7HDVF/Q0XGRDYBIHNgSZWfayj5kqlJD+3iu+/4ZQrKWuSO24AEBxSHDAXxuh
xc64LPUa8CW9rmQGzVRWExJ9EfYSEUsu/c1M+P9D1oCHIhgQA3C9Yi2YqkZ9LpDPsXJHF8mg3Zlz
2qpiEktZqjbXWejvckMV2G1st6H2PAwcE931FcaHtNoYSMXWLJz1G5xAwiL98lZDfFs83T+0q0D9
zehWFoztV1RrnMiUkwBhfKqyNBCR2mUwTt5gMOMdBppc62ZelXcggzT0LF7fNA/OHtxX+N+D4LE2
09AruVIJ+4D6/1AoRcjj4Jms3m3JCKSumbxSWKeYGafGDdbw7FyQ3uvTh207ZOs3rd6CBljjSAh7
qpRjBDWDRrG6Sb2c5egzhAixjQ/YHB01w9CyR8RVZT64mzoyOQJINTQOOMCAOIigsrv7l5t0FODz
WuKsSI+gc6tWAomG60frVmGgt22El5Go6plFeRGzBPX5+SJLxqwPF/fOXm6dfOXCR01KFuIWHt3g
3PhP8YBMyVglx7146gRQqModDvPlw1d1qRR1a2xmU+N3xtWzIqgYFNF5LZXyw7od4YEKeJBuYgMD
9LNhzCrQkZj0LiHW61VXINaXPn1vwXPWOfsiIFzf1mb5lw6BysC5vXb7haVAvNmSAyV61GALfYKQ
bK66ZPP2f5asHiiffJZfiNrm/JpJKQMhwGPzoLBbTD5N1C4lbBz3HHy7a/ZPqRaiwHfs4N3kX0JX
+6BRw5m+kmKe4KqrZ5F5sU5tusZXXJFwjFVWfCBqXkGdIa8Ya8T7QcAG9sH7g1CBOTuE+mg0U//H
Fy8JzBguqQPrbGu0bcUqhqfRF4DDORCZ6uuDII6DyEyZ474scO8ii1h/L2GA8xyg9GEpb1NpvGEj
xBByKoTvARLE3n+BXwfEcI+nt8Sg+BG5LM7OOhCPNmgnA4YsfsqETtUVRNOLr6SF38QKlfiqsGFo
UyS2pkNsY7sysmUlEavDqlwB7mjftngHgWFcL9kHA+HtdbslMIOMwWnuqrPE9frl4ZgH0QjvszEG
js3F3Nt91zORsBOkSspC3YrtQ1eZrgfMjXhHe/xIebEC9lzjhreo9/IVElvXqEaITTjZaAZ2uN31
wqH6pT0GuDUXH9QuOf6OPBESkyYtayV5PQBEKf5oY+usjMInIkUjfBNTaeIjBL/PVXqr80ivvKyo
VXbinSkRCSHpY5CFALLhPQvs0J/5ss2QurEf2nXbJmLW0y8QmhHdvWVYNr1ZBlZ5BVgitF7M8KRW
HY8MhNPE9kjfQaYVyWzH5PzVQSQKw1IZ+kK4WLGMVaDvwnCzLTryfqo3HpxwBQLacYxeB5DD6VTB
GY3Chc8KSF7TmrVW3JqD9sj5v+UWXNvUr7DVjMgdlfKvcZt0eE0aWyv6YoGdglDB9UNMwx9d1aR1
Bvzc8l7vLbn4px4jZhwZliru+YtM64sL0lcTjC6efyCtqSvwgJY2w9bQtkgUQoed96PqYMGR36S8
ksJSX7+pexvwkiO3jF85AacmrRnEaNgxJ3HEF8LvPg2BYpEU4IlvrRqefvpNfymQUTLkpsbYftf2
83CY90m6vXlF/dYqovoKIbnkGOECytHyvhly0uDPPhTLcyWvEN9lUeIQdE7c6SJREA67C9TMIjTc
IOPQjkgHH0A//q3Ybv49r6W8/LynC/CP6ZsUtG+izCoaA2COY0GqukkYVOZAZdmqJb/X8e+1Vi5H
DJEY9Q5HUvHAj+qOXkIC4vuMAhqGZ5Wa8bgpN3fulg9Ip1YIXlUaBvwlVGZSgL9v3ewbWljnZKRp
fsCGZKlSN/oCBJdLMZJqFAAqSYzf9Z4LK2b0FGpif73ATwg/OkJSjBpdMkHfb3IwSHFST/d+7w/V
kNGJT5izvhEsE8LZ9lAZosIHgqgIPK04ahfldUJPV4wLAkrgOHY+MBlVa2cMrp+LvkFHjJTKEGOm
f1CUHqeA7Dv13mxwUdKIqXQszBXE8+YROWnQWjSpA/ULoh+nlWKEY9K+2NW010RXNCOJ7TYvzbZV
yaSsSpPFdlpGJjFDknfaXENpJ0clxq8MEa2SDFe9rLuu6YPwknCrNHn1DDy5UH3fqmbKKEQSisPh
R8hshrTRV+kXpBGnL7KcIHOxMJ0Z5W77yXAc2oSsNvsktpy+NBBHuOP1yao8ggaWfpuiHDIQSOI6
j9fisjJAb6FLb0vW+wNql+iaUH4mHAB9SjiwIzQBtDIT8kplCKXQOqaGYSYSipHK0Hnehn2NIpME
HCZcqgk4W5OGPxAEBhyi05hb+UtyORMleY1Yphv9GCnpPe9Xn6tZIxajZu7sNqsa1GXs6/fq5LtW
QEJnjnQCbpwQt33bI+CTX2yBjESm8U+EdD7SUuPPLzMzm+eO35XRdR8c4O4swJ3j2Ke9nTXmGkzP
Swq1qc9VJ0JV6ScHj++lPqgG9BX7oP2fNS8ywKmMfC+tuexokxSUoQMtBO+y986aPH3qLofOVFcg
v1Esq2ghFeuwzzC6p14yG+Rkb5kZ/J25HgJBTf7kMEvcBIjahctJ/pTP06wIwTxBwt7Txrokfn+M
lnrW8I8L5oddIXsTfTESZHNJ7kA2CXn4Pky9QGCeio1xjYeGX+uggq1tmieUXDV1KjLmu6wUDG3n
qDtDT+vu0D4GQWOMQr333drBWDzECOKfo58QiyqkaC7CB3ncUZF8jfmyu5kFGkgF5rcgMb4BneDd
/i6HgNqdnFORF6fisj/BgK38vPEuABHdcUagYo1NQCP56i3vwqblFylEQ/X3EtFeafctaFJY4CXz
P6FMnIumHYX+8HZC6iHFDGsVDQMbpJ64KjexTj8BQk05WIzJIVInm4v1u2xh1QWNUZyLlyotN3Nh
O7CduGhZC3iIA01ChWvcnDfb5sz/ibTTv8oWaC84+i9tstNZeVHquD9kZxx9PsXv8Kpe0K2VZ5Fw
VQJhv8U6WRomwFtNtk3kEPfTYUPFpQoFmt5/KVxBpw5HOIAXJ1y3YTzw5ZCrTBhaX6zjVcONXH/t
+jCnAbjvdjKFG7YuUp5tmA5PSbt47JBpsSc/oM9Mm3yRhoAjIj4GmeP+qrEPo1dt6REYEc3CTD31
w9dXQ0n33a3AmQRMOBc22W0NsDso8Bjs31YS4l8sUQwzIMMYRoB4v4lTxq2xuxnSdaxP1r1zqH6C
quU+k06I9kLVtxepztX14okTFJ5b3XPeW6LKS98MK6/2gvgeZfemymPex21ew2bMQhDCSsjDgsl+
eMJrE3WBrBHddlJL/nawudxU6Tqv7OFKlZ/61ChlSBExKUyHtM+bbllyfGmoyeXsBljxciuS+FRQ
i4cT2meFUox4PYEX9y3QQk14tA4rOvXbllooB7hiXhVEIEMG5IWCEjbSkS9XPQQglmwgzTl+t/Z1
DdkyEXCo2We4QLA9uQ3C2JVwOz1jwJntm5MVpom/cgCc6dS3K+TbsPo9NKbcp4MsrZRko0rOFnXl
gPAeyoHAzyACUPPGJWS3RAN/+/rOR3SWMdFxlo05nXgmFW+fJE9kO3nfN1d4tDChcZUfUQ/FCY4o
3EcJLtp2rdpHLVZDDhppeyIxdYYznJoTIYXkd+U+V54Vxhy+JOa/tEkKEwIc8NllBYdeGVQ8E1Gv
tpkbEfhjVPXIOyhD2lt2SqDqqt5ML/RefFbsGhBHVDpol43oIqsG/l3xH5gxo4e4v8gAJvp4l7G7
9ax+cKMRAA8vOBuJ9v2Udz09zxiOdwn5KtgU0p5HQf3OK0z0z2Z27X5Jj+kSCl7ETtg9D/tnS0Bq
JLtAxkX69gq+xVHEajE0foud4TEXSL7KAo7S4tSoFOqlXlADOpyThqASSUtYQOX7IGfoquXUERfv
J7fvU++eAQz8SPsQWxba1//Z9zshaGzrBLao83XtvURe4R/8b93R5tC5M0hoDGBdvDKnY238AmVH
LJnYJWmsURLGGIK05ThROzBrsCUfjgdNz3/f+OG09LomsHOlqIgdIMRosAHoy3MUrQtcgcJrDhD0
9EMqq1PL4XdTXjSpwkLelF9bV0jtBHFS4sqFHCHcM8+w4kvnHnEgFR8dUt1KQS7SZNe6oiZ78RMd
NSft+/dSCJ7ZFmGzHDCmIw3+16FQcChoCWcsSfGrR8Bg06enXVmc5nHEBlvCspFtNPE7RmcPSDZP
RuqbQTlUgrhF+EeAJ4uVscdl18i9c4ERHh5ZN0IjGgO75V690jk1+ukHuCkBEmxa7gSNOYVRKYjH
bGVnWBbnqrpACI52x9DhiYHLNCUtokTFN70xNKeJ84HAXgobys+XeTK/ZxiKlmEbI1kIyfYxdB2N
jxPfScZLkpo08al2QNeg4xL6aEgPZikQ9deLMMp0gKpmfTGNbZoe8RTeLCKQVad9TmfICavoYP3b
A2fEVkFs0YxBx5Cd3DA+kkfSxjUDic5YpekmrwgTo8WYAkXO6MCN+rsdFW5pIPUPG3isnkqsiJ/9
bvVpUdUe+qYEFBdnrY6KE8rS1Bm8Hc2aP/7mut5kGJL95PwQf478vea/ZxgE4CF+PFQRJbGZXbq7
P+i0S94/+JnmJoDQqJ+p7LJzhSPF1zyt75mK6Yn75P8Xsa3RoLMCYe1bhNIooMH1gjNgBh8k3HcJ
GWW79GMEm6FBHq5eWGJBzOucsKT5j5SeZ9B5w2tv6XVVd15+HOxwHzDha9pNq/Qo1KER+chhIvW3
0oH3Eu04mtHia7tGShY7QiBhxFDyOD2AyGKcd64k/3F3RnlMDCzCMC/6fUN3zDMaAd+wVApnvn1Z
43lSaNDHvFg5du7QEQjnC747j6Xj5bb1h7d68OjKuKyg+PEGd+d8vsgXVuYh+cNKzwK+Gj0ES3RQ
PsL++lKYjn0ZWGOiwjfjmU8tBKM29OQgzlFp70DsOzfENVPQdehq1NziR72RZgePs5Iu+87vjiIx
ngpPrg7Ng6FXqwTDGKQGKAuw0upcTheAmu3LT5alYpkqaWDXLBZMkHVLUAgLVPWlMx/o054mnf1I
ria+TzJWpeHpsYMmMgS6eMNjxgqh6JqJfwA08wueNeN1i06I3cyfq4aANxfu+t/UrhtdBg0NJleo
GYngc4d7m5PPst3dowXTdjnBzbSjm1ge0y5DLuN2VI4K/yE5Apl7DJhDWSY12ie/s+FN39GBNMKf
D7Hr/Z+tIA/AYgwHK87/3opoSnHh3/cZOoLKgJrEXvGVy5WtaoO59HJ5MarndGA7dIT+QUKYdlJC
q9QrxyeRgCGzYfRtQOdNdk2nKRvc7Jg7q+cWsgrCQ4g9xjtteK2EcLfqWHugKjCSeFquP5/KE7fU
OcUSPfAA7/JCLO4tO7aHzppDa6mtVak4hagcft8Cxgkufx7BvfksnmarBuEGFruggoP2Pt0d92QT
5RmZ2pfObD8yP2yg7yy+PASpECLKbFpS7vWibbbsC32+cfbu51+41LxSLvNtFiOxyYIk6XfsVtR0
dmwsjkNMLgkuaPE/axOlOgZfUqcCe3ogNxJcCKQwbR6VDqF4iVKN9BdmOFUgTCVdqHpUz2RAOC9l
5LykG67YelDEbC/o886pSmbQryEaeo5QbB28H1+fk7J9slG7BpD5E/qpHzaOesIqnuX/QcV8uc3E
HzrZUZ4PuzQvXeKGWG3fwo0IzxKLjZo8o80IS87EnbcFzwL681pEl0BmEUzJW+UXZ8EKAHTofgbg
GznPq74tpgNIW5tjb4UBpT2P03sUEkatk1qDJGnN8OHV6APSltA+f+DNH0F8z0+Z/uibMyzUSnmB
BrdWsyZK8Jp0dg/TjAILEnxkMPSEy1bwhk+IUPx+42lqKD7oA4WB5hGKISgzr7J8sB0w22+5a2tX
dL3Bvq1nD9DKzREG4mbTtDvSA8USyuW/HH7TJKEPS3fRdLZwMWju7x7wpeQtVl+vlTFQkCmgWXs2
tUD+BMoBXeqhgjSVo6gAO0bA7EgmkTpcSClQGM9EIWlNL9HdSGvIvAiwsT5HfZkOhKQpOTxMY4X/
w8bBuqrWPI9PPWl+EUWmqZSS9EDMD0DmKzTpLKvRDRFdhQxk33hDtM7XTI9H6Y8PaKmERwXXQqmX
Oao3bunFxkWcWMf45bYQTqq0RvHHeYw/0EHxH1czuiiI7QwGREjI6cxfHhGehDIoSyg/gIm8J/qE
uP7XAejul9Au4WBb4aNAZnNV7rJu/WvPpmtf5HdV1gMgMFpK6n0bER3ZMtpMIagMaLbW5zOy8b4g
pevCP+qQ7+bwnRZNCiZzKh+JJiUQylp59UlC9rVebJlPs721oZ7gJZ/h/vCScuaq1S7jQFDzBRvu
1o9fmuImFBEbVRyRsw+apLbvLAhsndHntaaGza6jRD0PPbyGic5446MKLvc99gNMRLQ2/kjDsfrX
yf8pseOxsunOhF3zUsJkLRLnYlGXmr29G1LPdFW8YZDXNItuxtX1rKq0cI/6Wy68jvZcn9pQypds
uo7hsLx1C/Od4HVWbzwWGaMAYieuq2SqOWfX/SZuOuLFptIDIWDzzOa0NWcoAB3EGXVoKVA1MGOR
SaipIq5stQLJyHq9Ovmo+ynjYHAw8JWfNkqT/uGJ65YLMdmPchTCx+/cug0KD27iwaTeL0anNWAJ
6cdpY9Kg4OkhlxOKySa9nhNJ8y0BTtwXAnehbqzse2ePDrRkEEyiqAW5QWqsWocO4Jz53Wku/jPo
fjeg+roE8tuEb5hTD3iQ4LUyox3TpDw1DQBPBCl203MLq7L9mLgnU/Gwx3CVHUxFCqaOzrkRhQ5B
isiuhvB9HSP2r58IUdoBDUCy5pl75lV8rEZoCaWF776KbLNRAKnOPpZRE73yUwgP2AMrK9KUhblQ
8VLtaaoFCcwJeab3n3/XmktHTQsgY9W7E5hPVPu90C22heL+Z+yel6N0eXUyPLxwwIfsft30G83a
TLPW1Q1TsGtwIxx5u0CLN54OemQV6oEnOoa/B/93ewqjbFbcd0DsLRt5LrLo3pqWkRHEyv29zMEA
4xGquUUBlIZfRSrPE3ADzp9V2NdUrulduif7ynmrKjnEUmCZXxXMmbPdviNA3lans9Q5xhf6d0WL
G9/zfeSFKc7H3eSp2vZA33cJIfMH+mp21QhcJuSVTxqB1Xounxe7f4++Vq9uKSK9g5+2qqUpmVD3
cuAT8sZRs+2mwjXGdHar2nJGYIapo6PT4LS/BKFxMXvfDGMiqu3in2wnP/LXePc+1JraaVb4/XnH
7L7J8T3aDix4NyVM4rRbmY1L4D0xHGhZE8IJF/I0UwpAV99pjmxWQYx/wEc6E2851fRv3e1Ac5ed
AyW1bhDH68oj3u4pK8ld2gX/ymGOxaQsJhSVDxdioEjVE+t0I1iPmsdlN14xHixo+chKgXQGl0VO
R2qTAdIT/8YCo2Zou9MEXIqo9joBSRmbnSOHJ9rfVNupCD0GF7mZtMGLm2PVjcPJ26NUprjWOV/C
85ry9GhZyJX+LFS/5pCIgJFkTH9M/VLhXaxQ+sFwcHq01LEATRp/UB/ufFASAxlf1xsCUic0NQqe
Go/4DQFfTgAI3fEwg8Z5d6Wl3cWTEfWoh9vX1W0TdaYxz7pN0VO/X0SPcJSEXVMw/E8b839v3dYI
iZmlyfhIhzndQ8DNX8SVfIAzTOclvbiBav0BqmWGRYgUr7UTXW/ER1ym5QEytPOhX+Kz/UAgNpg7
hxpY2ZzvGu9wqTrhNC+KmvD3Oj1XkuuTRwDC6ee9SnhcVIeq4F/RUQXBrn+ejpym0N67DDq8ofgg
wDjWk4JZ3yx+phaktr9mvsw2lHRf35hXj939j59Pg8q7kcRCwwJcfPVm6TnIsak23LFoK9PiZ9Da
81oFlU0hoa/GmTjmTzUDobOU/3JimgTsgjUypfFh00zG5xhS/I9dMbiOHm/WdQrQqiFNn8+7me3L
z8FO3UuHQE+35N9Jy1PfBqMLiJH5g53Z/EGfRKkK/dme/kN/HjIgbDSzvbUr9Fx3CtVPpFZaFfVT
wq52dUhlfUnlUwoKrhAPvuYQTEGwqxelZN224KAci5s4wseey5zh5GH6ThSZhWGwoHSPi+UyXYHC
+h/Hsp/Syv+83obuewTxVNFFJUbo5MHwu/GlAzJE2qJlP7L+2fg2beRX0szq7mP5taP3eagcWN12
r623wBaysCeZtmcxV9z/87stV36Kv4AbMsFnskcd7zkbytCIqkvwStzLoACUuGW7zq4brE5fTYH7
3LYA+WA62biWN4Pp8JHqvRp5aCXepY4OtykS4avBycDowoBFABRhOxhuoTy2XKY2rQKTcSTo8KeA
6bkjnqkCs6SFG+ALoyIJRTdWDT0OUrGclJSthB2JmDZv/cB0K6fnZQKbRbto5ZcP/W+rT7uXzQcN
c+ok5T9Lps99+6w1pHjHvb1Tu8JairDXjEjZ21979BO+R/AIryHKYeCEX/s271HyKfwwI+axMRkE
p2ZMP6/1lE7ANJjndXgnD3FUir/J+a3jfIR/wT0jVXzBXmRdkwDE45Gh30y9jlh+YfHALGoxTSrp
g7tZTkYGz0mmZaTlGxJNgp41MTT9qx2Fa3d+GZGqIjXrcofZggXhGQTLoBaN8Z2pT8ZmOqsLTAds
H5HY8FSuGLbb5gN4USQqLpemeWvpVrf1fMLxxHNLkWsO/7ZAH2At/nY93OGIVU/D0m2cVDkvqU1v
Jy4oOE7QMPiyWWpUDahSUzkUgkteSNl+pmh1U0tq4UGHYUwJqtz0nzKA7VXbaRsPr/6/9hZ1LwRP
UN3+aGEo8R3oSe9IZngQzdH7FsYEUNkjQdWYlDsV1EddM+yhn2spbWEgTtmm0Sq0479D+qf3n1AI
+o2ZVLtiWCktQzGzkFdRsaPPosKkWuk0xHjhFkiUMy1WXN27CDofDtfUnSeTW140WS5iWF3AOwFr
M20cO5qVfcnwHWPXBd8jzTlDPGDCsDAPgFGcPiYL+uRaVU44/BiN+agdRtL0CLICINspL/mrZHI5
qIMNnbgKCkP7kePOnbQd9OB6LUGx2tN1O68rBXcJCXwsZICCVDM0Qgf9dkolZB+dSfae/bU7D/Jk
69zPwcjkn45oOX3tstHm3dtBFbRAanyY2WWPlNvWQeFdGA2iL9qdGxRikz/jd7DDdmRr88ou12ql
Icq0uR76Lpi6Y5lXG/hM7uWQF3oMnG954CaR1DfRapyc0hRSTDDv3cg9YHCMacM8L8n1cC0nwXD8
Y47NNWeKoyJ9rKGHiWmbszYrPYXNtePbzBPxzuwqeC9M6cjNQDDDktWMszf0ygtxkRo/hrZEU7XU
9sMuV7lftR4+6uNvnSaabVtK1wQFONn+r//BpDMFk/ucmV2xNe4SiQW/xCdN8puzFptci5VoLe2U
+/PQNhvRVaCAgor2Ip2sppxN7haGz6cxYh3qSMNgXxY5j+UpGhJTqOQRW2oenYSCbbYH0T878biw
N0i6liIr+39WdaJydOAXy768tDrj82rRO2NjNXxTFWq/jdoK5VBq36k/s8nGoo51ZK5kBNqyCj7i
nhEdGxY1I3rtvCU1WpeGtULyR/2FN/hqnM93Okk5MU44fOazoB8EP80UqgFFC0+YIvJrA0YrYdQx
5eaY+Ih4Iiumv32gbF0BAoAnU1JF/WxZP6CLnb8yafRH8gq/51KkeIxA5in8Y4MCE6L6Qdcut11J
cgA9uUu0ejpBOUq2+FYW3QpPjwLkzJnngrqEo9kWilF4o5rYO5UpnIhIkINQE+n6Yu1HCHSB0ft3
N7W4kTIc+HAZ1E1FQ5mzwz3fU0Vq0UBAbqmjn4HUUsj3A4f0+1y6P8602fJRIxNpGw438sxeXktM
bns0i/JLTufvFFeQ6OIlIPbqulanKjDg6Jb35Ehas+kZKfbdX0SGh3kAloAMLf2kRD+i2NN8Zn0I
eYVrmIQ9mnVg/Lc7x4unjM79bgIHZTvfjhKi0K0nCf5/RGtRTFCf538ZfbyDZcdCdpNjY8H7ivqP
qKXhawIBCVpA8ZZye7DNOrd/aWq7UEtrxurWovY9YVr+4j/0cMirHIuK4VCxY/tnwXZzB+pkOCKO
SJHwKdet7B+LLcuea7kwcrxSAc9gHKcZd7FG93DleyWMUH02Sn5fsiFxq20FSAKKKLplqN6OKy73
0qZLNDz7rlLKdMooIJJk3DLfT4b9wlnasrVJymxrVVBeHNwNTKQS59j5gnjV0bk5qGLN3paJ56b7
amTvnbudfxdrXdNuvbSsR9VQs1i5NqKWYo+0BV5S5295N+S/Ph8bXeHTlAhyBTKq6MZHIttZGWES
gC6e8wk8+Po90o5nvewJ3NyEmUNc+MeZygFzeh6pQ84MS+GuJQX7h2GAArWzc6pDUVjtgz7EYelI
up9bKm7C7OmaPOBouJC68lp702QhjnP+s67T21FPOEbM8s4bZKPLHLjhX7w0TmxmPUyIGH8MLulC
e/ZxxnxdQtkB4QIW1DYXcgIxzy/MNDzx6t6+lk0/sqKj03yUWLLemnRJoeS2/GNsitjN6iiWGZ2t
9rWYsCP5tX3yrri/Eap6k3ml9sg0YMKJJSgBzCzukUnt+NvC0/ADRla4gY9YVEqCNaRleOlv7kRW
79BxzIDdwcQCHPJL1/4s7Jac90QxdRbYXMt7zm18iOIr5f2c4rMJpqBpmC7eAyzVf91G8D5CpF8T
gVrHmXEWt+aCXK48Ieolsa5aywZbK7USLlXq7AC4g6Hn968infiSo9gmipNQWpYifdZJZzW+yv84
IZMsCSTMPvdLPulkp4RhovUYRqpQ+VteD96iLaGXFcX1Jd32w1QI0gQV8VKPspFkLT6rH6mhFxpe
RxX0hXGvR+0s6Xv2L1K0lo+jOD4tMTo+2wu1YnsWhQvUgc1ntgSmdevMSPl7Z1SqOliiWdNN7NMH
fa6zSRwt3JI/U74tnVgVp6/5RZvZllRmTCHd5x56r9nN/MpYSZhtzpvGkl8VSr8MV04Xcw+IBtr5
omwAKnW3y7w3xFgsUR73JrstyaDSAZGj5W5cLvjUsnK8wMWtflPUAUdVNXYZYW4FKRa+4+prgbaa
AkKx2fAaR7nwmLSgCUzH0RLHglYmtrJsIASAJxLKtL7Vc9qXDuMerfMNY2LYYVF02MNM2Gkas9uh
pstjqfVgLA7QZFfhXo0Y4K4Ga/1QPbVO1THNmJnv6TbS4BIpO5N8ykf2MbMicQBxCsjBDPzVCtku
OtLw5mvEand4eO8Ml5y4qaejU3mSR8uyrhxqxTTwE8vaDpFzeQeCpq4EpyCbHX1acbpsZ/7p/IqV
t2mEmIkYLHgeF8ylk/olU+mBFfkyGR/ga+ayItE1f/WxneRhOeBUhk8mXM8Qe9WqvOeaT76Sb39q
61vgcDQq5j/8nzIJO58dEiYqm+TWWT8OpPR7Zh6FacgaoMq4ie2X+/ixVB58zbSuiklOmJlpO845
QmY46wADmKPRF72WDI3EgYXFbZFuuzm8y8I2KTGuRUM2Xmmopu6QC/UuBQBhpKrsKcEtc0REiwN/
ttpfTnae0COL2FMcc/ad0okb22ccMy/5cqB9LqjUf04h7n0sLnamhFJy43cWJ5Pd+/qk3iO6OdRX
f29u8Rhj2rGGEAmac2sNrROzgHgIucaERP/6uEEzjRIs37Jpuwj7wK9VeVplSv5N8hIvvNfmHndI
hNiMterLOCJkHxUVr9hADLMvp1ugjfAJooAcSDvaxAx8FyzNwqDXshk7ZfPaFsnsjC8M4VAg0jZG
gE8VvSPQvykNA35YODxbNZ00dz3WDG4LPphDEBmKY2n3VUfY/uLc9G1w6xigWD2pQeC407NH4soo
dtlxn//WrZR+srG9Id9g3wILnh+vsTRdfYk0PyFkxs4Rq03EJSTNh3M8y111Jl7Nk6ueVVCaTWsr
e6yEOLGUcwNugxj36BN5X33rdGCD7vZyHh0bodEhvq5LvfaNDFxa5LO9PX4btcWoGAYTCQY/YA3o
JmHa2cTZBoKKcCiOyD8W7U7VuJB7UluLboDyOCmoNIrX1MrY6SY7bi1vAPvqL6o5YXvhpFqAhQz6
yA4Ycdtc3vmsu1d1PUiRgMv3fYjYJ5+TpTrYGn2sSQ/tjGj5+pNvvfR2NTqK0Sc2dUUzn+emynUq
CajG2l69SrnBNUfuisuSgn+Ac2vmLnZNY+jx7+575SVvPw1yh+KshqlVY5T6BBUZMekst92WAPGL
aTspP3YUQaL1gVa/4PkQevagDZr41QErB4ylKF030UfIJoNs0JvMdDJaUN+I53sspO11lJkKsJHO
rZFNkWkJ0IsF04WSrVs93pJsMpJOsgEYHWyoYD41TbOM9u1f6lRDGgfDnxwnzMEpN9ormXPawr0J
eIeQDJs7wQhPP7k9MTLSRV9p0xw8kJMuRh04YjV932RT978z4aHDusDIUlmgLJYX4381JNZOP9wH
Shr+TxtMwZXKHVbNyDEt85y70S7ABn4QkpYbvatjS0owzla87yXAvYQGEqyy2RIl60ztQt9buT0d
DKMk0+H/k4ANLFwxq5AOM113yevqmuXcOvPWMnxOIUmNUuC8xHf/ffXAwjJoWi9gPlth+bt38JK1
40xy6U7XHRPlZCjCalGssxLDrWC2n8v3fQoz5ZE+2ZkdPGs9YbLkpoxUmGX3eJXkr6y/4yl4s+jd
513pEj/Qk8gqJpa8DA0XmmQ/vD+2aSWR3KiEjHqDHGTSMqM5V3y/zeSsJelN5iZXhJYrxy1tx/EG
52ziftaZllaBjRVruPA8Quju9dHLM4PoDjOizwKCnF2Pjb7gXL+otl9rGmVbwU9YVhh1Jei+nOyT
JS3mvaQVQ9xXXPw569g0kW03YmvJqBpUl4ULZXxDHfsOOxUfwRLAk9D0bD6lQtvIzx3LrUPVh119
N5QeYaAnnusaJ5WLZn03zU8yHGOv4W3o2kO+m10zJZq5xacayc018o7DUibRXgTHMOmzsz5kNIaD
/NsaZaA1P5jueDEXZ/Me5q5LShND5GsYJ+7OOK2XhSw322Y9iN9ZmQxsDE7S9cuodY5hSB5eMS+r
TdgR9e0aPm1WEJ6gwxbQKBuSGkqQ/B6iYeT1w/w/igUEiM65eISLjx+sT2IiXG7ByIiBKR0bxxkd
0d6000pLhm1XPKjrttY/f9SqlKvXy6AxusI3echc6WBRlk9tL6Z7KWapskWStQ216jnsILuAQyRc
NX7iAwc91FE5yuIkTjl+4RtguccfO7KOeP2iyy9BoyXzQc1Gf9ozZ4IjuDsqdnKu96cXvVPSkFgu
jPlq7meGk0LpkdAaW1z89IOp0SNy6nhZGwLNXe8V5T++TO/QypNqL+ZDklWZ3BstZw4FGwxo5J1D
0uJJAymLaMMF4sAlvv0WshSCdyz2zXwrKy+8TGmvUhJ25/YLDnK8sIFdnSvDwfXeSMAfvoXW98E+
AMQIFi/hWQddvZcW1yticeKJrtTwN1G59dIlgnO5V26tsgmjZE7znxk/k7jIolxFJAGE5IuX4AR1
GlarexE4AoJ0lfJHKx94cMY09h+f7TWCyOXY8lZnf+2Q65MslMcwu7SSc0lnuLRYDGmmz6Dd9OsH
5KOiHMhS58GURm1+K6RYC14h6R4Io+3r4dwjG4p+MBTvRyaKy6nO/LFn4og0N8OR1xz69kWYeJdW
QG/MlTSgNLlFjTWyYF7239NUUZ3X8dKksfeq/Yq0lQAtDPNJjCdx+ysjc80VvBK8uDe05pEtOJ3v
7i7ak2g8KbwYFL2lntMogtkwRjdmXoDs5I+CvPdh/1gCXUdyrScl9wSU29CyoLRVQqAvCi20ntak
MTEPa98KMBExcuJUSL89y7sEMKmk6ep3yFkmfDTRmf9Oh7aKndhAKnc5ftzzKzaG+FlsPkBKCzOI
OFHf7+FL/pL0rWwTkdIzoVehxWj6v1uFhXxFyzRKXbJc6fYJbjO2EsXLiGf9r/PXD+1XRjn4j3/w
4uZrufYyywFSW26qklZ/c7fJ+2DdDHLuPY78Y1hKbSKtDIKuisxTTBDzzGIqVX2LAfGaQ0nQSQnB
IiXJXyhLZ9LBj7AsjJG4df4TcuioWppFGF91krOTUwRWyjZ+gIxc+GF1NmSx6YgVKed1ONhxB/1u
e+qzuECGS/3TGS5dB+ER/h27xR63Rf3AwnYT6Ocf2UOu0eqmf6VMZKpdYE8w0qf9wrOyJ0lzQ/Yb
vOpVhanAgSo9EVb7gU9IBK/4cSc+Js1Szd2Rsvc5wqMFGL6aJmuXja6grbCKNSrxGbHJK8ygxSjb
k+Vii6LLheJ+kO1jBp5l/veDou4g5MfwyX6yGAk6s136wWPmIQ5vXBGD9JfH2BujB/qjuBuCu6iR
h5/jcNnb77Mmo0Ah0oELBJ+EorJlpSUdBelyU3DsVLqx3fXhnhOEtey9n5tLbLHAWrGIYDin6sX2
4TvgukQzNQc4QqJ6FlUdhLH62/T5dpvBGzCGKgRzvBvSxNb276AzDV+BfDL6UczxL9gegSA6LpBD
ohKKzrmrUzESH6r5f6bxwpeDDEQEqk4v+yybKFoZz2GyEOpXUSfHd5HaullpLSA69sTr3kMCB0Wz
kpX317dGLRLH22F2oov7pcwOAUpAxQ4Y9MmqMoV0yS0PalcIY/nO1Jpmjr6IOXigk7304oNVVw8D
TFcfPYdnDpnG8wUJtH/iLyUkNWlXo3xeVG3kFb958Gdr2b4Kwa1EWb/plfGhmWPNRhG/Laeyu9fW
T4iZwAzQv3uwTGvmGW60ZE6XqVRzMeq2+W3eCx/mrQE6dOPp+/qwdDIlrwIfYDKI+19kL+Wf3EEv
FiIppRrPxE+UwJseFXOXJpRF2GOd9rNik1S05pSFY/YURL6y/LLzwXQAM4bkQK7pfBQclxewyMRD
hz7Sgbc5Sqs2u30TuyOD4yMqA0GWuPzcJ6NNEXSzJUZEqU1i517q0Zb3olyMrHU2KSmXvlaQ4OKs
GNOZpzhSldfVLQYepyxkaz28v8oQsF/2VAuk27rA6yCkUIbHnqhPA50hv2yErySER9oIBUKvjXh1
Hgg9KJxiWcl4HWvcolvNNa9mRoOc5W2IPaLlylaenlOTiDYaOP2MW8pUrEO7W8odwGDi7mqBZFeE
gjtWtX9sKtvJQG1NY+V+kLyz/wesdLnAVpEc0i5X4Msm6q0OeprqCdHVQ+vDr6PNYUtbJw1q54Jx
sE74JEgPijboBHeyf8pE7niYBGjt6wTmj5rKBe5UB1eYqJ3n9sMKrkJs3Uo5Njd/lOhbnALGQLM7
RaZQTw0199GzQ6KzLb1bJtm7POA2HeWuf13ejOyYEfEqeky2x5Ljik4eLGs+NAtvINaFO0qEdQgO
+E7NIl8tCFZZtjXFoT0jys0vDFgs9n4wrsM3nNbnnqNR6+iyANmM98Y/iNemOqQFlW4x3Algj8ic
tBKGBFZSHr2OSBV786Qet83siasXHTv0zokl6rCJZHpAPT7GAaoSz/nCiGxDyCpfgmEFRvgcvy6u
Ve48zxo93HW8i6qX3VQl1z1r6Sen9S/QW2MoFFPYBl6gdEBff7tYN3VclPkGdzsgms/AZMflNa+6
4Xs3mFbvVK9g9kCVVQgeSikO8RJDOKQrtgWsnt66a/mWaeE4G0RalEeg8VE8C71ZvXCxclufk0Uk
TbmAbbu1sx6sHxxKHoBJOHF823yoxjio8NWsWGqVSeikpPO95H3OrUt0XrRt9lW8nfssOu5nsD3B
dtAqMDrwrhySkwQsLcsxYiWCfZvu76pRsB1weZWwyVxUMIVXl1uWm91FLDGh6fjMqEG/o/B87oZQ
Gjvg8mAe3qSHTir+PmuemurWvFr4C+E3/7CsX0H/p+yLhG9m4EfTY60Iiz9P+FykVO4+5neLlsmx
RjvT1PUAEQ6mMkvZgj6uHes05twHT6dz8QbVABQ83MFzLAxJZju+oR43QjVZ7QmkBJpU1HShhhlU
ajgq9upCSplD6agCC8Yr2+B0fP/fs5UKSi0CSjR1A32QSvmZrNQ9482qeRPnChcmG6BujT+1ctAW
vUJkwbU+hj7ZCtI8GLPS0fqoEZDR6wFE0hCLY8QqmWN8SjlSJTYIPUGyl9AgS0SO49kxbTA/bWgd
b+S1ab31dONrtyDdk0LcncnQmX0xCQoT2hx3SHECUbUBnuBG/axtksPwJsLTXMc0QsKQGDQWz5wU
yNjGw4XpQQHGouDoZv8OSkr/1/RsXdCeJfQtOFt8NUbb279nK39cJOCWrDP6/zJOeMkvkkubbJJh
Z/NZupjW5gEIlA7Ei1eATTCZkzfaPQPHr3h9V61QEElFaNYvvdAaSHv6shsBZd8BuTRuxf6IlBaa
4mPjBk5XpoM26lkyZpdDNs2015z2aQpbOx+Dv1YvOtIjEVrF/Pe/x0arImneBKvB7kHugZGlBGFO
5xHNvLWbYajOHni+77h/wwEZWoHDDPkH5lZ88BOf1y254PDwJEq0r9b+hZnq13w50pXRRkWWShwy
bv9EOjuyUNZ8ISKNVhOVEdLU0g9LNH/DteH/EFjJ2SxoEeaSdYRXikebq4GKyYlSDh0qd8XDtUmo
Am7ES3dW54sOfqxdC0+dYndsBQSOQ0MklbLpVgFAIQN+0vwKWh5LzuFql+i1TIqMs79I9wpTMRay
hyrvh56CiLRYzilBI20gTxRsOMcIPBz6mUzxNuKARFrogvNW79fhORf4aIosjkTVP9SoZSEXbE6K
JqEDAOiuD+eaRigimBBY+IXKeYhsV1we1TLzmkCLiXwVm0yH5TUVDzv3W0BJZmgOU9dzZp7ns9AG
auZVUw08wujBMdKj/VvO0CinPAjclbubGbJyqEiiLXUUTR9YaaogMCK36RA4NuAGfudjmDufXx9V
vMumrRSa7lQsp7yFGV3MmeM9NQ7HY/W3rfdMHBn2QTPcqKlUZJ/yOr0hyCUCSAh70GbMSwZxB+Eb
Aj+1h0BjUHUKKJvTmVGj2vlCPLQG5K1GhnFNdAJKb6LaCaiLLnjy4fvdiiwjfMo0Uv007kd4Xizv
4PlVSxkRkoqJSNO/aqDQFOawR4poERfDU1FAaZs2iZCRLgTMpaDNKtV1YiZJ8DSLPQFjG0/PshCC
tpArYuClSEk/WPXWZHk6aYNJ8NX8O3jEZTAd60riQsSUw06TkTBIoWZMANi1lJULEcphNtcj1KkH
WnwDRanBSZsAlYzr323E3cEzjLMLfzx6Fh90NcmRwoRLoQMR0fWTSDuRSSmZ+1fLvHyveNlvEEQl
2dPJWTUUei3W6CuK0Llu8ODSHphXQFoPlPBXcXDOX62sI6Z3+4EICo1wk1z+fk/T2OzSzpts0Lvr
R2PW9Yh3tnq44otczt5Z+rR+gBtYgOZh0F9yc7H77SmAggN3GGBNhKuqDe5/N5SrUNsoZri7LZrC
EEvpduf9iTTFTG57bqSLyznGYd1pfChQT1XXEIeXNVeRNk6mUgGXt7ne9jiBWQ4OeKAuzJZqiUcQ
ikyGIxI6mi/q5BVO4emjs7r1MLdMOBnQlsUb51DRT6ljN39xXCyMynex55bkfVLpK5vaeOE1YZZ5
/cwkXiNZN1gkHiKa5azM5U+wdPzFvrT0OQqrDZNnRor49/V2qdAoWCWxxLCOofohMSt2EO7/81Ow
4rb5w91OtxwoLKcc/EUxTpDQOirTdMXgyk2H469+xm7Na4UplQOlY99D4CjJUTOEP19eAsyyr3B6
CnN1kn08jG+8XK0nrr01hbtjrBnmbv4W40B54F1Ceok98lyOezmy465+HYaHC9u8bbujQPydCDri
MCHfh/AKRJ9GbF/n6UVRdwHY7TvYky1ixRKIPE67GFeQ67DzQ4z8fmbTtuVnFzjRjpqIqUVa2ZeP
jwu0IeI4/QUDLt4h+ltS3FOeVysj/wLQ1Xf1iQuL9tsMhgNmdvYn9IZSoeFb713CJJc6LbZuRTM3
dn2jQlwSKowyKJihgJJKqtwTPoYQzSuEYUnqzzipwOxOPxxtXSyTNY6nQkcWQMFuVf8jHXtWPcbG
fuVG55B0zv9KXQcpmLVX8tGI3X/oqnp+pbuOtDPM2LMt2c2J6i8t73zvIRDE/p/qIyS6JAmf8WsP
wUHytX+1mVUPmKPfE4T8+biHm3yGV9YfjKmmctcTAwtdx+ibUwrtJOuvAbuxmUS0CSvL22Gn7x12
EXtQpurf+p+4CuCmpfY2C0qAlxc5FDcTA7ONx/BxlJLaocS38v44hPQS3LT0q9PQWfXnPP8aBXn6
FOEvkkToILRbymvcGhAuRTMylPtRIKbvW4OvZKSJmHCubOooikuFT0WRJxk5/YREF3YomZnAyFog
yAudVGJ0PwZBLSUWxGUC9NTEG6RjMFNVoCMfygUn5HcKgZUTQB4OEWTQeU+EQ/zCT2S+IFGgxwZT
w2Ig2/T6/HH8mnBgwFSaC4fOZ4blwbp5MODxF6woVX28esb/9uuHuRJQzTCh+DpMgq599TB/b31K
tb64chnI5x53+DD0zfl0AxRdCfCZlSpZ0klN2oihkHaJgOzT9jB5ej8wW3EaMIcYwPrlr7eiPPEI
jqqsbZEZVpxwxiJL4Fa1mZGsVfgaVp9864Jt+5g6gJfJQW1EDOxuUwdDMAQFEspVSmxpILgE1arh
l/iGlD29ptAiBeJSevQpTf0CCK/n4etQljrey5YwPFqXhgMUBL9hQ6Uok/SoDtgfXh7cG3psVA8C
6G+36GQqhmHtfx1aSOdekFVeIrcp1ovVQjiT5hvrA4QYW5I/OqTqz3RaTj0syow9NBdVTs8kSTY9
C4npchzEHYU9xF+3w4gjiN53OeUAhK3KzeZtTqu5rC8ntuI0UsGVn/0ic8t/EVv/4omz55FcGYFg
g32Xt+xuZGkjnOlA5uYDoqxK0V3jB5Vt6tOx1YShAw9yR/oCjpKWt58ul6s73qeKmJl3tvk3B5rg
7o/vh9TvU+9/ZRsw8MomzybPpI29fmr3iflghSCV+vAwU/aHEvjc3n0q/0YrMuTz9t+0ZKPoc6AK
079pOziR+YLYMdAIkuerFAU5EBjD1OaAB8Qfz1oStB85jHO0PtOV0RZLs4/l1WVM1FZxiv5j4zth
wplCs4QbVYq2GcuhUNUGJwTmr+VqcDN9FeDN82emLLQwifpQYyZmghXyLo2YjeaS7RoHiF2SHzBw
nQalBbuyBqKzIy1HhbDTlceaD1L6UqEKPa3NDK5YWj7jU/d72FJwcpmK1ill1tUsZ3T6rQ7Jqy3D
Nd5zXrrUXv7EEVjzVYvLfT5T/VwFg8ljDY0bYxpLwwn2km/ps9sXiSQCyxMd1P2NGaiyXNuDZKKe
9UgdrHk0Pe6doYkV4x59v8jyHUbZUzFdJWStIX0x2HeIzQ1wcNibrlp+g8x9U03LtZy93t4Y6uFT
zIKENMxw07c2IZMq/jBKYI0y4UjL1VcH6E9QZRCLc4rvU0yurF6FVeGnHQzp13Vjm+09ia9xmgJI
vKYUXISjKWidSKHsDlLyRRHDI+3ApCwb5ZOfrRzuJGqhLjQCARlTVDuW3uxcqfJdd2RkcEMxxaOA
YohrgvheWWnGHmliW4yQsF9QT6XT2gJgza6xe1E7aEdjrWAS28/gE5arnkpnRlhEGYkOtP3JOnNl
olKqWrbAo+NvzsasmZhtu2pYQv2N9ygir5NKimi+Wy8sowcjgtB9rf306IrreO8hW/WJ2gF1wlI8
TrpjvgYqhEQ5/M8rsr6QHXRwceOtk32359AJvcOlZAw0JFYnFqCfW9rK20KvWKau83MxLOerpJI9
1b4qzCQ2Gg3u24laBYTNeYqxxNPb9bZzD/SuEKdlM+nxbWj1SpFUpoZTl6Es2GucDQ3jyU4Ulmxw
VjR9OUOcLtJuIUrDw7YfAbgLFb/DIa5+RzCWOzF+7vn/n1pG/bHf+1/fmDS/i7RwRxbJ2zaZsTTA
GQ5wEYP0N/RnEx2nxSdIczSWqJGtVccFkCKLneCMrXFOJ+JA0GdVnlxUlJ1fDNoF2c6gS1DHIrUl
MqHB9K6jow9fSfPGyKvGADcrJy3q3xBUPqg/ZRZf20EKxUuEm6P7iz3+X/osyjQZwjFsrpbenMvn
Vv3gXBtEE7kUWs0O1V0XjyK+0ibBnJm4Nxk2K6g2fJUwdKCTyYC0gKULTKh09J6Q3knkY/geeW1A
WLXufhe+Id0KKQO66dIzhX+o8g4ouMhP3szmRXo7V9wFdZbOBb8yXo8I7LxSjng7giaD03BwSCZ9
jYBAf5WkaI52esp88lcKAGat8/s9i6ZpoxBZ7cgXzbuPnLHl3XKUAKi03t9ta85IULNTQvtndy4l
reR8bwKvBze5V6Rok8DkQQtjRgUJLiS0Wgz48NbJZwEC8JeiHec2/+7FJznl+GxCnqBhQOxSjVl3
LFwGR6SGLJGNzNJgr2xGl5yxpKjftvuIJIAyo3SMqfyjlaPzLnEGyXrZ2TGtao68xF2bvCNsRljE
SBkq3XDq/DZawVuLsw+7ieKrSIYCojQzB+n9qOmxIl7jv/4FNBVz+REOhmqCwwtRiT82CsiLL60/
HhG0zGCL94AES248jVdlaieRyk+6PeFAXvDSejkXZiaUrX8kEQQ0HpNaKapubxFfQiMCyT+v6/M/
mn5t3qZ6omm1FF7BcR6FQaJo8G/rlOlbk+mHthLcABx/riqoA2LxUBT7rVgegeQnNMAdmo4u+xmx
q9dYq6D/QkSwOExmox3SUliSD7kJcdqGN+/zaqlwyUfdjFZdURdLuGsWwvHRzOheYjR4g/HGVwXL
UovgezuhzAbuVWNQRt11gX+1CeMwl86K1dRgiEOpNvZnmhqVoCNcT7RFnB1vT9/M8Sr26a+spK6s
xCJjlz8vwspfhv1ILBjoLVtxpXpqZ5zf9RU8rJ8BG5hf0setuA5fKFGbXQ0j8sfsC4AKnZJrPxd1
ea9uvstEKaoUBvs+5BMzq6wdOFafNkJhYj7FRFvc4puU18SiRczaBKscOxcVwCnxFlDnj8eoggkj
IK0CcFlZC1rHOdL6qQRMJePN8cTBF4110rSKQJVoaOTMlo4R9spFtOG0JbChPA5cuP08WOSCBYf6
+VGnDmYWlKP3ZdLXcvq42GBo/5qcSeYdJshbmlPJKKDn1DON354H1v7ib4NJjUFEqticrdWANa2n
YCzsqPrRwbS4CoEpHyCf5+U6iVGmzCI6hChnVUPAebfnI8BSEat/qX1zTEnncCohj+v0Xxj+NmTQ
xmEwLOpjbRakI7rF7GARbLzw2GIdSAoXAW9RhWZoQIgL63T1VUzu6be/HbZD6iktTtjoY2hZ4I1S
WlqWsyCBy+eW+d1QDyqMTJ6T6mleWikhbIHBCxUSCevCQdSDyoPkuI/QxUT0IAbYS7dzmOxMqG5l
4D6W/KYixf/r8xn4UWYHB3tcFe9242WiEodT0p37Edw4WcyA8vAFHAIURuWRKv34FUd8CNDy/R0n
rx6G26i9VRWhqpnN6nRboqClImFzDncvqkDsSr9EQIbcZVn3aF+pwMMcY8SurPpdWsaM39JqyEwj
o9uw7SvVtmz3Kp3bOG9eJHwDIv80jD+DUB0NrbvUVVk+0VgNK8iU309whuQIQTjsgkltOSOL7Wah
BKNP+wdhezj+bxK3wnSCoyjyOANySmaqVfppq7iypDYpM8Z308ERZGNlAK3BLq2iQwgtOxqJ52lX
x+4vouZsa7oYZy5AnGpr34qLOZQ4WKjmNUoereo51o7//dNfElJVSGzu3hI+SYqoA6lk3QYbmbTd
qUZ32+Dy8ufXEK+q3kEu0NO4urI8/RPT8CF+N/LBjMQa9keqcoWJqRF0Tp1KeoFz/+6J/LXMpr9n
NCV4a8QebpB25hBd6KHKjlBwuNb233UOeSdgOKO2UvliPmCMWAGJZKqnYcqMm+CpPrfRFw57fV8x
8ZePVwl/J8gsct57UcZspkgOZ8Fz2WAfuIlJ1KJdeRhQSlnwUHMLhmJ+G2qULeZoZy382Mes/lWg
Pkcyz84IPRnxal02Ftg0fxpgEiLrFWtQ4dCKAGlR4qdMcLEYwHwKdBONTh1INhlSNgKEt7d5CEIi
jtvgmJnQaKBd0gJw3sswISmAYvNoVtkzOcj27KqqvBhVKJhF8AN+4Tb0Ck94HRViPAlbDEjtj9jN
Rz5OlI/J9LzUc1G3ktEb1JHogsFuMdp6ULPwTPTGo7j7zEwteVPScecE3N/jEiUyOR3Qhf6KgRhO
wkpaCjTkd0w1sw3gO+yoiFdczLo5Ckj86bp04Ik9QtZ62GVz6kip3ca3O9K2CLJ4aKfUopZFcgFU
NLDMxRuawql9ZB092TftuXgB9MkN3TOhXcpN+RuWkMoijSCLjPQdh2ndUBMNkIesE0QKRwHs2PwQ
VD1wTHfXWhB52qzjuDx6z5RVAJ8bvMt5K0WR07bU1rvzqVsTuenuraDyPQxtM0fcue6bEj2gfXnh
RC44IETrfYKhZYG81/tOWsQRxYtf88P9mG9QoM/9P80w9RvdA7ZghYL9k4wH8jmm788mTBC2yVcV
YRY+Wyv8kRkTeU5i0Uz3qB4wixePcSvvyuEptyzrKyc0z1oU3tHfajYAhYUZIGkGw3RQ4/S3JQwr
2tk6u+aT3MU8ExnWVtqBS45ABwBjN4Au8XvptJYrN7oYuMK/LmZHXXevEdsVPFO4kfyqWa5zKTwb
8maV0lkAGv65XZJFSvpaeZZl87ZWXgblMZ8/ijLQJdusPM6zek2aSLU8v2yCpjpfg5ZsPiJK3kfF
BNMF1D6ME7/T07zGB24ikzokK+54GZPhAeHzhiOKnIyXbTBvnKGOUkOoFc1Ry2q4KWjnBGeUDurb
/JXXF0aKOOBy5sOJ9kmltpfHx4suAOt61pNUshWtJe7bkpD/HiSJDT8cLTKvxdJFNbtbJAeudfoY
0hH78cn+i9pKtPAbj0dXhgo6RU1BgWiyFH4cSqEH3KzC3QK0PeVckETi5RBdz84dxnlJE92E1XrD
yc6d2Pmy4MqlyqwXfKTIVCJSFH+aHdWgby5LblPtCxPnh7uBeOYS2P8eSKvWIPXdN/Y8Te5rNkp0
LTvkAwYswthTHMx8yfxt36MUpviLqJzmmB17bKzZ+3iOXZ5iHCtW6TzwXn43uJSbZkvcYvA5zUBy
0Jz6uilO0SBVfjoi5g58fd741BoXJa/TKvra+7dWtwCcVQhUGEIKPoLLTcQl6e3HSaaOy771RYV+
OUuJ7TJVZI2Msd5A8HnsZBaLoNyFHlNKYhjVg/xHXHPgj1uE2Xj79ITAXnNLQq9AF2vLOrVH9BtQ
ltYeLgU5Wx9JcoEShjERwwWxMPnVVueRhXVE95eRzOX3yjXzq1hSkXKziZ8gvDexJfDy2mAmWrSP
uO9iMDIqxT2B6cQrb5EsAgcHfegZY3piaKEdlVDNqLMA/mC0lOdd2EF1L9b08ubVm+0NxuQF6+cK
Z2p7bPd9CaO85fL6QS4civuGd4pHRagR8qwUezE91726f8VjcXZrZIYtJ3MmvuSP7VAmUdDvqbCj
qyEo5bVB9ubGb1qaxlKbqAiaJB35FoxYSWezljgKfZ7gLN+E9dIN9iDB+d/WIDIXFYwmRLBqzaEL
RTL8YgwjIU111jJAhjM8I06hFEHNRHO3txdfJINW/wRVtH0kmpfiNRzzaECi/eIpPYh9oPRfjUV7
8MMm3qh+3h6GcuIE9HzafwpN46MGYn7hEORlykxFjjxqJj/KIvpN5ej9FHWIOFStaabZSYp0qk7L
XRAtEhYoQRuy3EtPKXgydVG4CiZ8NcGAjOl5YwIxma2XpqddZj52CwO5TzP5K5oas6fx2pI73J+4
necGK6ABmOUJXJtmS65WK1ZxiBJH+fEwfoN19nGcSi7M37GKtTYpsJ6NQ+D/Kv+uSTh88RcQNiBl
XtyihBaP0ZS6Yp7Icts76MZZ2guttvdBfNZ/D6b7n9tLkIadgrOz52/ZtRZ6gf+4UtGnamCASX5V
nAPhPK/7WnOv4YbNd+qENXi5JauxIAX5FGAvKzQxrw2r1PpbrD0X/eLegxOwTwMTYGSaSKZjvbIv
lAtgvyTMkOWSTdwzs2nQ4RR7ZUwKhHzygnMeKiYD0/GdOf2MQNmleo2INBV3Dp/jdawtB6VrhDIF
uWRwuZiTxF97HwPKYj0qt8Ip9NEfIVqCJ7ytbFHMJhIfQnLLjLgCwtxnQcVhELEzbg4H2r3TwChO
ocg5B+e8hbsM7SW3qX5F0uXfRYmlfvwnoqVkm9o89d31icTE7SlsIJta14exLzTcudboXZLdP6gn
F4HbbeA9XKWn2zkGoM0MY+JFIOvL499SfbwlscFJ5ODeo+sPPMn9DG2fQutkEGVy/O7jgDSrVNzw
S+9PV5TgoHc8GF8oVylexr07SIWxLllnkqrn6TJ3ChNPrWeTW167dC8SQzYxbfknvUITHFM2RW3B
S1QlG3VIGbHwCCdBsZoF4PyBSIRbPQjWRkmSW9V/3vRN5R2oq9kxiRAe9cvi178q/PKfk4UZH2O3
5d+3sAMb8x+q+5ROmFvEK1u3udiTy4pVcGqPxG5ekolvqsgjiCCM3tuYqncDl1gWWrAZyOE9Fwab
tKmdXuULiCasSn6FH89AvChHQ+S0aTsJweJvU+faSlML2eDLLilE6anfGpqb31lw4hPK5eva5Ka6
ZM6a9dEWpDiudCNOPbtI1w7CYKjpAhKvltYW+oxJeR3fbY87TLtzzAL2mo5qts2XFpHdzl/6VVxw
HjDLplgOnd8fcRfHvQPJg5xcxVkVBmArOVfGSgLhAOfY6WOkxt3hgwtKaTMo9NzWLohVdCgomg5F
610asUbjdu2mEMrRCvo4PkluN4UoYaSK9mUDp3+LTw1qzBCuCk9//MddhWg36f1a7q/xPO5iWE0d
lMLdnebV/E10sPoePljjXE/aDzarFSOII2H++eCOaMofELbhkClyx0FuwxI282JyEYz6yxBY1HTK
qA/pY1zzlfSIAX5TtUBwNoQheDje+h9z0LXochuHPTSviG6gB6AV15Ixz3GAP6r6+G44Q2sx74fK
RrjcckxkmwsSshK4dR319MkSk2DF0n2E9fF1k2GBANUZqRXxRcMQSxMsmiSLL25EmwueFOWkavEJ
DFgOzK+N9bHJR53PLsuvoASdDgERr19atQlYCEGs+WRJmyj14s6kp6twW2/lDvA9Aw2yH4JjzX1H
2ey8WHshpKlNmfr4IRNzTVv4k+qDoZupd2dH5yiKO0zjcXNNj5xrEQdwgUUL5sxGCUEy5NMStPoL
25RuCvi5K2hEK/IhvJlw3b0NSOEAjk3beEAYZGFUTPDePa4B4Jk5QfaWZFWW3lMpnBgW7KqmcV1p
hrVCoDZynEUVgPeyXiJ6c2JORwp6b/JLj9IrGAIUAUzXl8ZMnlI9swZaTZePvuLllkYxI/GXjh66
30mmr0xP7MdGM/pzekJjT/dC213hVBVK+XflJJuzC8g1TW5GpXnsLcXhXzktIBYw6VWDGataRfC1
mvxxG/zd9Wr4MlQGSF4cVt8Dss/3fBrvie0kdETYXNR6K+/YoyMXeQkkUcNxPqwPMPR3SxH6AR0P
5pQn8PnwUHjzWnWbAHQDcsS9cwt9RpIRGHQjVE7lemuw5IG7PeSCHE4rRK89eJYCV2mvUUbBlxyY
5KcIs+JFL1iVUUyfauJ1TiDNLyqT4girz+IbNQ4M+hCJSkNymVRiBrKxYDohztLzK+pURfYEqY/k
8wKQBYM6oB2mcJO4geMxuRWVkbBgcB6UEZZFWIcobQtosPXmY76vCk0HA3+RSvhjBP2a2ThrcsY4
mtFGqFNDqp7sSzhe8GTjIvJ7/miKn1z520YYLVV4s+HqgvFl663z4rxO5hTPeMHLX6TuSRiUhfdB
vis9nOdte+x4Pa6E//X+wLfIxe6sxy/pF1nwqTTJ0jkjRMrH2InIdOB6mNJJdTEB1zelVRXCljVG
mG3kcc13ZEVgC6CXG6I/Hjp9wJQPY7eCW6C0W6Esj0pQvNGkE1uKw8KfoOthF9wXytkmoatJc5wn
sW4wKT23Fy0yKJvzt2jrIthEqskP7NTA0gBLm1sFo1RHOt0edTLPXFeMrqhs4eV2BB5LB62Jq5um
BG3o4M1pTq1iZY/4Hopwh9WiI28kBzgzZOZ+2blGPMbzXw4yRvDrJgSjjaLEcNYTAg/nOYpWkqAf
gP+4Smch0Tmuk7awKiksDhdoQSVVcKFW1jmePMzxypkNDdXxpCRkyHodxWIWmyeGLokoh/irMFdS
5kv1yMO7ssOZOSfU3RnicZ4EnDHWkvpPVurfpk2rTKu+ysfQkUr73egQtrsDKTU49QZ75tr4WcE9
pXJTVGOknmnLmt1iPcX9+tYUgSeFzft8xmRtlnhzl0oQ/qF0eYaa0iiuV5ngBMR1pWH93hLWqqYe
JJUg2oDZwJeUpUJvi1v9M+CY/1YLaWHkd0G2khVujgBv5UcGrIgPKhP/9qTCrROZFv/VPQxobMzv
Hvr/XGHNcITGfR6GGLmyA2FBe+7a3Z4s836BJpDepgrLafDp0TTdfwpvkzK5y6N9kpzRSLnV1CTW
cYHG//fy9U08BvOlYsvxU/oh8aENo0c6tDjBSnSOxUHza7OmWHPatkNqxfWXuHeXiwwNAmgv2Rsq
zycqYbF8ujznoK4ARE1zlzVCOrVDgLxl1oRDssJEfJcOPTGrjqPybC0EYlQ7fyr37oLVY9kcz7RA
bgLj94f3uwsV4YkaBe370yrObpkqShgY7tZ6ycRhESRiTmrEFxTzlvOJA9eQcPyPDOGGP1f6Avwk
bLRG08XHT3hIsMzXAce8h6q6x1/NWN7dVREO3nnpbzZNKgxPvxzcdWoGMg7OhHoouN0u3WI7LuxB
WP/HBY2438ggNGWh4NdF84ndVEtqPEbjf7MmDrhYsNcQH4YY3Xztotcuv8zeHyytNblsGhIswURQ
eID8KCESskQaEhKq/eXUQB9vR884sbbQDogbX98OUSy+SmaPGEZiT0lfOWXuP3Y7e9JFJhQT/FWP
+kcnq3y60BwfuC3SgYaMS74Cha0ppY2ak2BI/oMYvOS8jt95AsGEjAuxPVftOI3yI3hNDu/93CDZ
YarJqJa97YGwyYZ8qORXlJ83CA86L6O9wM4vXOn8reWNUtB2fYhfUu05nQx70mgHZrcU5bfWdHxC
fJIFndUxsIxUa9MzfA2+eAz9a+NiFuhTcjNrT1XOqDuDt8CxnfM1R+H4F/eDpELVF+TJTw6FcuxC
C04fX5V0cm0d/n2/qsYxFPDIIMHSPa+afh2TgsOLKYiH5oI2NyyZGKmbKlns13qmGPtRiqGzHFEV
LTH0q0JJTwTBFjMtxwDb0Lgm5n+lKiCoWQkodhV5hMxT4f5R4nIHL7DOaOIpdKUavT3ZnSUnQtgP
GOxXxeu8mQPsOJ70mOwsEZEVN4VwbeNK5DF8vM7WGnJZhpRz6fTPTkHmFW5Rwiz2BBimwYbB4kxm
ijSFmIr/PDTlzuk2/WhVh4egTAU4lwVoW7KXVkBd3Km+CqZEX05z/8A7Tn6Vc02pkA1/DrpdgpUu
6JJxz86+e6x20Yu6KHRtDGLUJ7bL59g4BK4QjECzBb/wV8Asnn+/xMbeuaAZiX3yA+KYTRCQIVOY
Fo7aLmGWnKMPzu9+SYe/g1dAWsQUUob6D1/T3SNtNE+FzU8ZGPcEhuwRl0eP8B6NS2b4w2PgrOz6
a+ydGRAwPDNwIhW8M9UPqYkIxCsuReJxHd8GecK3j1omeGtvel2u5jzYHwAEpKRHkGLp27csC3F4
iYMdYlsRshA7zajxNsfF1GvJWx1FXa/qTlpmisIDc+kGJc5Ai/IP9epc1bSW7rJcMrRWPHJJYULh
3SfFZHa+HJFWU1LYr/mZ0JHAAik8YUnol9Cp3HnoDQhVgvOmtN1gGzmDtxmVg8c/LhjjO0gXm8Nl
GT7Crwr5l9q8xC1TclO1sDr79O+77s43TfXjK3tomrXwFbHBfhJX0yMBBf39MadJuBVRRQAK6c7u
Z1vEzNb6nWFHFqDVoo/oZQ7yQvmxuO6pVZPuUlIcLOfy2/BXCFpsVhY6GmTJNQtiNMVqp6h5wUkH
ZP+/yH46AAnHnxkxYD39mFSertWErpZdCs1L/uhc4VVrSJ1WROYAGXgXrv7fUn8VEr4UmwA1XSDn
KhoJ1tCR5kPi3hNGPZ/bTYVUiDXhizviG1XvqcR2ECr2IN3rTdmG3Mh8J8kca+ycTqwJF5GZntBJ
nT14CLVm5flj2w6NCiUnZdeaofdyAHxqWrgQK99yXKqBZ1QcsZBwvfM28CwpLkxtXk/orHsAhrNG
RBS1X7IIiGpC9a4EcTuZm39gtREERoAOKei98JUde0afrkDDWigu764bCUhYXx4Jdb2KOlXOq9nv
WJK0AvrgukfGb7h9ZhPTlO2XMn+AH9TgCRUqQDAJ7CJcbGjxNoS9w6dChRCDMHzJQss5uovETMi6
Cv/59insljPViZlrsEN3o6Z5L8NsK5B5gY39Tcq5k9SiX7uSoQjEwtS7RtcWQuX31/ELr56+j8Sw
NOvkQ3GtqoWYTQ94Le3IxBUv6vfttPeDladPyOB+Z0npEimMewfIKv3AFXrysTIx7NaKV663Jnbn
MuYIlSHbynzWrsSPw/P+GXcU7yxcRXk6pfpjMAE9hFIxtMcTHKa8bEKFeuvVJTNJIQ60Mh6At7Iz
NrBX25uv4aHA37AHdFCx0fNF3SUUpPM4rBfcFwr6F7+3TBBN3qUG0p3mcaZFjz2VBSQWqjivSstF
C4WdULuL7vgAwIkiomWvmQnJsnb+A1WMvsYSrjaha6TENqbHYEeVkCPa6LxaU6l6DcT2rqz4thSC
Fb8dKBiXiIjVVFp7iM8z/X3fg1X8y3xH7I8DiC1017br77NugD53hj8REPpBG6SC6ZhxbIHEVVVz
ktekr/b1uOibZjQWJC/HbctKcLMQtNANNPwns0uNJfLpyb/sjpnd1sSsp/RZTRdEXx9aFIoj2bF6
U9HaIuSrnaxauMOGoRBUq673G81CxBZYRvBVK/BTfgkJaWXWbuih4y/jWlJXzPKvBV+Mabw68WqR
pw9nhhZm0kbHa70DVRrOPRZKE73zd02UCRGWCr0O3KWvCaH37ZrgxejofJWWUCy1aFSPemxEbo/0
oMwLBL8U7rv77ummVg3zZZtQaLwHQKwWPDsT9i7i5Oyj5l1AtvPoFoJP9GqdvTUa7ASYV4BFI8G/
f7UbCFbG1WCOfIM5SsC1iRshKPbzvQRm1vjQFcWLtIMcx/qA/7in88c+9OQ4g2/3nBDzPEanFKNr
4ZHpWHnt6OvzKoKLwjwntkjRvIgFVyuXQ12znxl3w99z/dHoh6MWWo4cM4xO2KP+rQo/aHKsd0fc
A1rrYk6SDb75+T3zd0QQqDQ5pjE1jCW55LwNvxXBLh0okEBv7ErWdZMrVcQnNvfr/Ys9oPB+Zkbe
00IG1tFKtKMT6YICBiE43whdEZFiczmL1QN7pUK8dddL/ayyVPM3NDP81ZtEkYc0nU8gKgmCGjRp
Nrt5Z8Qnm605/JhPTmJIoX9c8J/qrMoxw0W/MT6MyNMMpETrCdJn1PC8DWoBQgUxQJCKcG+386D0
KHhYBMxVKk4CjBwgnsRG1fUsOZ9d90T5Dc32wLeTF02R8GwbxsWjCV5JueZcbMFLGlpD7+fm8gcU
R8sZlQzQfTH0gzOOxxGddOoLYbCnueKY6EK+lMsE9YmV+5nHmEu6qfWLW1r9JbWw18YQ228s/n4K
D1ZhB9XoTFjzaP1VBP0OmjLRRFndlKr92hCLXXIS73117uyddt01HhPjpCKjJKAV0hF2L093Zx/7
jcOVVITiWJ5lJ19+boT9f3sV6WNQeNpIn+TJfvgMofPjclL4YV5DIVkKo4CO9PajVocdrEC8DlPt
VYijfQR6OMDXU4iQOE6BOEQ1yAs3B1eYe2vKJRtbKbl+AtPUerFJoU4yU63h/oANOkZ505XLxVas
SzTfgxhX94b2HR5kc/CX163hi42e/HNoJFRWNOHC5yqrI1Q13ceXoi+VpKfSVbAqaBiDSyTEZ6Nu
nBkB2bm36Av8FSvYSHrrv1uDGElLa/YzQlzepqMUFAMJ4Rxu23fJsCPKWyOVT6GlH9Oz6y24fORq
Sk/6+9ETQVl0VpAxO8IDnzYdj14T2XPNRihZJz5vrVhKXszZvftmXvec7TvCoT7VtScecxJA66sr
Zpm0yCDgmjetG0K1KTJdn8Qk4Ljs4A5GZxm4+OvIJSABVoASt18MDl6p9cTjJuxLKpJw2+lBlSl5
2oe3equudrzeUQnrUqa+FILgUdbSUHo7PxqC14CxTexF0Gu00lQCk+Dl+GW72yBALbDsSfiCI+RM
TazGLS7RnHfkdT844CDL5ZCM0G3UoIkP49g4m3aAwvwdjPBB+DuZVa3y6srzT1Xd/C/r2LQre5xz
2yeL+3PxmPhck++Si5whppp3UyMRIB+l4FK/MlHyJUAhm6WZRA24Q+Uqb4fnfagHWz1X0wl4cdwB
z+UiQQxRD2o80ISWhkVE2qx2ipjDTkIPkmGtxRwPDfGpD/Ux2IknPgcGSV2foma8aqpmKuow3iKt
Hhy8f6UWrro0OE36W2f6My+7DVjjKjvaPk4Tw+hl6c2FqYf0b9B3Wd4ZyEiiaqWs4Y2Fw2xH3Hhb
8ep8l9ucYNzb82D4kySzDE7AysVIY+/6C2hOMqdKHuPZpH6JJYA0/XJpDU5ZkBrconv3uf9zhXly
6wASsRCMAY4xkGNY0TrXUm4WVhn1l4GnQXwH+2ewQuVAJks78vOzb27hav6MoonqOjT5B4Hd5XJW
/6w9wwSVyy+GCafGbDfbjXqp7QxkwJX9BSkME7QpWjHydJSxq7v8oNw7HQ9E5r2mNi1jDJxRESwa
pTWlgqfmWCnHjcfIhzPF7f+pWr6rMbQDn6Wkg575CQo4o8byKehbHdfZpbrKCqL9KhIiklHxpZVt
9ZiS1UIF+tOZ5KLsrzpaPKbq0r6Zh3JShoz3HmV6Zrkc8h5unaMh1mnSbz11fmKPK61nX9imdydt
GCKAOhYZmGxDLxCNvlzF6TbUIIBiCuhsFuzFT5bLg0AqfTmssuMSzVrnW9HsFgcYPT97I03wbkts
kUhFBIJbk3ibPVbXP10v29OxByQqQ0tmatIQPwHINuOnv99b44AmCTrnb9aEJ2JnqIH/7A2RRyAA
gi7moLoeMD+OAKZqZmVu7iWUjzMGajvE64drA0UDPJgcIa6PI4SFmwcZVo9GFBrChvBFtQmm7Gzs
PBip9D5p6aVIwe5eIWjAm9bXx3MjlHRZt+vE0W4HsbhOm9HvTtAQ4CLe5YRqdVnEbufRdF8VlVX6
bmcp8t3Q3G9eTSHrbTU/ejUoB/ObY9Sm6vAziZwQGQYj3kVHBvZYyaj7gZOLDnriXJHcgp/3a+77
ZXgVIBDyvOh0H4u+2N17zhLBtDCyIn0HQY5A/OZglLOeGI22mbW9MKoxia6ue15X6wQm9bD5oWp5
RErN2QK9HczUTuN/sfuBTBwYmX4ZOeYJUL8s9pGC3puyVctDYaOIoPt6lWrYBaIh4po890OV8Nni
DLOkDebTQmJclJV1a6BlcZLAZAedCbbxWGFeH6aNOPNQlTSKCy2AZicUIf4O7tVVXMmoSEdmL8d1
/p4wR/37lM5GoIQ5hMltjnksPinmUQb4ZRpUlUcKHwkgmHR91xJS5e6uLZeQIdE/UEiU4yRe7hUh
qtmvxyesj7/1PAwwUuFjt31CEZ8fi+BeaTlm6DN033/9+qLaWXz3scpT5r4RMwUF0d9DUy4TDx41
HN4YQddgeb9ucHWvrCQmQZ9QcKwxSfYwxLVjK8KriJ16tRNpL4fMhSYVC8pS6HwlTFFLOwymk2i0
9UqRinPk8bIFQSqY3NX1qZPJpSJD6RL/pPwrgRRRFgUKaS83vXwsHcJUTWYLPWaCS/DqH68ghLeh
WNJKpDj0JKOx+5zVM8A7oIqmJPfmjttcfVsDt01gSsa2/cvMVnmwoMNHkoz2/ScvNbMaQbqWz5lE
uFWIT5XrJCSUk8RMjO7Tz7ZZwZfdot39SWmL0BTO9cnJtonIEg5HVbmZqID/HnxiiQbA6JWVRsxi
UzabJcaQt5TeFb3JudBC8mbGFjKBFX4HFz/ZsUNBFdoponm2LBjA/ROShqJwqmRnkh2QVpzReLUf
Wa+v9TkDKWyl+/udNvcv8s51MAMZOxUK4v05Zt96QY0Eqgau8r67DMhPBxtL3COr7WQRN2RxYV5c
f9FzbBebIcBIIq4k2bMsX8akOtHahGQtdI/8svvqdx/roHmd09e3OFPjZYQXaYZpgkWuDn+8Hn1f
q8Fiw8fxem/TgEjcEmixeVAKYdawmTH3xSJl/N+0hl7LbGYtsWMIT/zqnU2mC1IffnudCdBKaKLE
ym+Mh1tYWiBRG8pUQwSsX8KdLTCFeOEC1Atxy8n6avJirnysltnh3PdUejEZEuDXLxqvXChkFRsB
4nvsxwn2NkK/saG1MV1qW4h8SJoUjuOe++RhmOIHHH2D/CGfYjcu+V15cwew46UUCyYZw9rl3zry
Uuz4+UnBqE6epYvJEPg4zElMGjkTX7q6a+MhBdBR0Rn+o2TEXnhPr74XYaE83d8JbmKWXCUIvxYF
2vf5pX3yrw0ZkpI4+bhtVr4LIXG5lh4T+K4uKN+AMfcnyckEhjaFqNfOcgqKz1afxJLzK0/hiqzM
4XC8rXfC0hjUomRGt+iEymHW79htOkc/zr3QucV3OSVhOYJvsqOgBtnkU9t7QvJA4Neu5mbvIJPB
aEjjllICn+6HdpxK5nwPzT4Jlzl+XuvUnW60NYEPd32vVB1NGGhvhW3JX2Q9X/Sef+bN6tl750ve
WjHQfg+bz2wrleIt6U30zmLFwDfneYeU8CL27x0R7XgkY1fwrwLHw/xiB9v2DCwoeQvnYV9dbqSR
nCxPmcKol5W4ZND9WimZYd/x9Z5xEGqxas8BPQ8i8WlmgPPVL+GQ2ACDhzyAZ39kZX5uphtDRU3c
49ElaF50c9gq69ygsM1CgoCy7N2F0iOOz3a/60Ztuda6ajq2XFUOkUB/YEJ/44fR9YBd9BV/xubt
EpDPOyPp69CV8L3uf8mf6bctAxcomXBQdBtUdCDwCEwvG+BVHU7no2Vk6CFboXjdhAUjSJlzlwYI
5IKx1P0r19IAqsYQ873gWE6orbQ3MOuDXOrHAslecOKA3yY+j0Vuiqk6WaVDK7/WrCPFJz62P9r0
IopyApd8SAO3XaHPjSjjAzFkOZBhrls4+mCaGaQJlXjyv69RgPFNEd/0k5SJFWaYvj1UEwvVbVUa
Xt7Qj7rg5xWunO8eU1AMrdtrJRI1YKcT7qKlom44nWg1q/xFP1JtPayihVdW0T+40e9X6FM+5KJQ
7vpm/iRq8/iPDgz39y/5HrOQSVLm268dK7Ls3Yo5xFBFGipLz7DOxIXDwn42LRtR1kwFUN+JIvI0
7ae68jGFpUjWRqSVBST28im1ND/qoCUuPY9Vclgix6G0E6+wYd8dh8naAhUSBWlr1tr/E9YZgG7q
cb20iEfJTHxYynKXScd0NCNIj7LJRotyoHO2ObPX5OzQFU+b+hMoDEMZ1dtNPTmWNP3uxmTG+E1r
AEwrrxDlkbGm3bq82geDBdgyqf3y5348LMdYhpoUv0kH59q4sK4CfLgFRXRKHUGEGcoqwBwv6LXv
sJsGAGISv8UQzOUXjHxrQlKx6XYKl6CaoIHQIhVFSWcj5ht35I2e+nD1xlBwCCmVujoQabYmk+bL
xZPQL+dbnT86iWxs28EpHJr/M8W6kJnJQwDObaqOgNfTpG6p4YKMRkazWNzlFbzorhY9mAzwmCUI
RD1NPfJ7vJwJtoWuEu0NKGVyJ6ZIC0yzTzdNzpoOiwz8lR47oFFvywjzXXXw9HvBboALHFsbHkgP
gG+NDNx0NmiUTfFinc7mQG9657Zot/kOr7lb7Ek9ca0TcRftS3D3pfug7GWR8DH1apo5EfYCdIjC
YaMh0hsFEYBJIo6oPRZFIqe2W0aaYW+IvxYHmmVGoIEU1NHAcDkK3/eAJwvK0G6Id0OBR4bsw83E
MCFQGlwdC0WA8v4HpNNwJyIvCkMpizIn0NdE+pA1DnVpKyDwCswaj8ukkfMb/09r5xuPpkiCcIGb
Xv+eU/0k1VXYlPKDF+mKHMDaHPQeipGmdYD0LN/ZTNvsE2XTXeZU6XDI343x7fGXIA4X6ysLyO9+
ptIwYp4mjCIgK1PVqyTP5PbvBzYLt7CkISj8w6C4TO8aOyOZ8vL66oM8JECBJcwdesUtlNYoddQy
to77Z9UdBaiaCqVF4p/Uk2EqoKzN46vi1iyp3gKXEEcaogdEGcOR1gEy5iOoZm2XjQW0yiPQyyxd
SlFTq7Y0oKjmIPl+PczPH/QeB7rhMQZd9/Kn6Ud0GqdEW31cfKuHGMM3tmoy5+m7KqqrbsdPR8X5
4qbbeZe3BMrE7MCEFtZtmoin3orA/pC2L/aIV9J6zxRfyR1AtMwc6p4nY6HnFXps2Az/QzmvcLKM
Ft9rwrVK2fSEVfMiT0jHFrQZptf7hD9Nj9u/BYKTZ+nQInpJRQm3C3f5q8r5gHL8yscV/Kac43ce
me+lg2W0EeWnRSqqpvXH7YjMMjZFU2V3vgq6GEnPTT8RWWdhme+rsAoyfMjKWxD9xMSP0Qumye39
smRdcDYW+Hi39/UeZZKT4fn3rXcRD1GBh3UlZefO02xUpJHrHr3u4TcKjtXZDVvX903bOOvD8jRV
0orhWpTgWAQZsDqBDXNoKSEPtoTa51C/Rrn8cBfEqcXBLmd4v9bRcXqETsoWkfLBbiWzSyUD3py4
uUBIfJZwDLrekDF5PnBjNLn6rEPsDVEiG7sKa9MRiZQCX26eJvhc1EMSrtQsh/0LPCUfZ1pHgtFi
MzdQlIW6pTijtAVT5rPPpoMmvxataMCApm1eowGkb210t3KyA25mpH57zolSmXqxhZTLkmii1plp
bpHasvbgzdDzgxdXSvXayC83yxnZpU6Z+XhBKpMtHbH5JdjqsXc0H0JjWiGrSKgsJ1wI0SuCUOUB
MohIkZvITMxrNZzVwAOSMID4Ss3G6kjKKYqSUFfuOsr/PtcYw3BJWOrSc/AmfTRetvQMpvCSPrDe
vDy7MLXKgZnGmwbUK2cSkhyobH6LzLLGRfjF+cTRec1D1ZSmUORx8F/FNVS0nRBszEI9a++pbwaZ
wl3z7BqoZ0bTSYopKUeEO0nffOo37uxupOZA10UDoZMaSgQywrlEOL8rKM9wThIHUzwykovwF5eg
HZ8BdSU6uo2VSnrE5plQ6NL7nO+ayGQ4N5alc+sn2V1VDv5z7fTuFXgkwCJBrcgLHMgJfU7VeTjZ
Eby+gQ9wIyHIcDoPxvNDbG+AEkxCINtEaDOKaSHwe2WN7IiUezHUbBVHOPldOKxeZ9GGNS1nRG4w
C4/kuXQ1EZh3sIL43vA7Ny34JJgIOFoLj+Z88t4y99EER07PP9e4cO/5lkaT6fCzQHIr7L5BtKOK
JEi3Ts3TFwrzcP+5T6z1OPV+BPb8xtk0QmyF/e8Y4b6l5cn93giPGu9fWTbYVb1BXERdLPCvVoXP
RIrCwKRl0y9e+3WZHmh/EHi8dbEQJPpHe7nrXlUvOk2asyw83Ol+xmLzZaEIJdyG5lckUB9cRSud
sqM2CxnESjpJceRwxurhdVHQzMu1XEuAF7pmd1tzeeNIDYPiTL6e62Kgonakp+6OupvqiujSmACt
jgCmNDixLHZ2/GM9uG3gTjIaeZ4yvZGjIdIJfw4kzB1D1GpTnAFe4t+BVWsOOphzxXH+fHpXhPQ+
bNLKnOX5S0/hhPRzYV+EbKx+Moaw7ngSsUgbUoGNTFDpWOSMhZ7LU6ov4PewhIlX+kKxTJdKCu+z
o/bbpL+crRdrXQ8uwkixJ5pPevGd7PkjEoLrp1Db6sHSz4UiPfmq1ghGhgcT/ihr4btNCQD0+hgf
36jdzAhACmg/mJLoW9/jHvZIngyi2uVxS0oKS4dnB9s4kbj+D7KHqxTCzKKfI0INY51JhJkr6+zy
r2qKMd5+7XLVEQ0K4VYsDIvcp94fIpQVLN58zAGazvJop1zB/lewm40mZ6g1Lju+gcGaxbCQ1jkc
vDxviahV7BEwyHpB7GVKTL+osB37LjR/YiOeMBNvvZb0q0GYqIA5fw5+Iom5G0d8kNAPOfnDOLah
we35gw+sTCUTM9/P0VK6o5D6ctKo6YJJgs1DX8SoMwx5AH9z3Fy5PL74bU5S3UYvoNA54FT42TVk
XnYMoTMkg+EdJwNBWL1MISFwshj267pOPheP1TElZ4pfRYlMDX0s667i5d73BNuZGqInLF4DmKZv
LoSJIXNCVzZpzD81JMR6bxUB3Ah97e9oXI0kfwjL7TMg5y4TWVbvJ9rpzzGj/VBMvSwqCDrvfYdP
IWtYFqPXLIrLQlErFzMdVJctyQoiwKh8Iz3yCbO66SEt03Bo7ubJPJ70b5cIwbv6BeHYMqD1xoDU
4mgw1Ai3zQzG/V2/ynZKR4ik6jqOY1SO75pU1NnAjEpQeC70tMtpL6fZJo8epH/aGAvWlvNoIchh
9M2OOpKycCIrd/1wXxlmSbPAeGz/8v40M2h56UYQRE3pDgiHebbe8S4+CXtmyljje1LtpfQRBs35
jC/7SftkmiT6bcHPORXh+6qnWROIMwhALfX9VjFJKnqAcJs94ZTW/YyEF9Pu+WA6JNia3BSNdWtv
X8QFcwtGyqyG1og+2Aj0pM36maHlwkiUs6V15Aj/tD5dR1jigiDagoWnjrp6INVY4GAHeQHjkLC3
cMxnF/zlD//Qqk9BKIsa5SvEbw65AJit6FifqGeWaQw75vrouEAgDjxpSuJ93nC5larAEPqZfKv8
VTTdH1IkTPrqHWMs4o4MCbIv7ErQxpg6nuHBAeJ41bYXKmabxPw/9XaXrUcILIDeSN/0/YQTSFuf
Rdti9KYBE7dIOq3qcKkffiHVPvpELODfYPUXQsTUbz5Nsm6mSU15Jlu+sXhGyVZgNWL/8amVKyPO
xgGtlnHvzOPXmIKtZEyknT51PaV+TX0p3K/MuI9FJ6TrAS/uftFnQBSObYxahQX1UbDJnbQQx1Pk
YwZrAYjDbH7nvnl3idXvGcnIxctggdvfOKaojmzI+XRxoZk/L83HTyzGEZTZNRv/5IF8Eu2ab1nm
zdcHB3b9LspjIIZ1HQ6TiLraUAzWOvzdqVOfVBVZr59rTMNmO6g+fE3NaufGTZ7nFr94rGjUPW51
pgGBfJ8BFSc2fJZaVpkZU1RDFlq/Uojecc9ELtTue5ZB0C96Q21Cpcjf900QTgq8/k70SAOC5BxN
JEk4uH7RMHDpT8KpKtn/J+mVFmfHZk33pK3h0vaGMO3tLB7yf1JDU+9TTcTNktcSdPk+YuhooXqE
EyO5iOB4ZloGKQD38XI0jMy4E0vHea6PvNFIYGq7b5e4Hc0S6Zwhp146cKE7wOqeKkC+Rn/OzbU+
mmgkQtiZmFjXXQmf3OJhul8AODMkEc1LuZ6qKeMTOuEYbaYTUbOrvxeKvmrKfd8vQGoxj19LWxgX
kzX9q4Fo+UoQ/po5QxqjIy4D1gpXKSR4gOlMzqwOOrEd56lstijCeXoCjbyZkESoWfAskoWiDld1
fbW99EEJU/ycJ4rapNyoUn0/qiK913GsQNOA+OA1YWP+Mxq2uc29qqD0p8sxZ+rkcejGdIBioyqt
JfwdYlSpsz1h/Qg5dI+P/qucYldM/ZwDxNxMqj94IrddIVNAUejz3SjZhNxNBdOqaNm6LrnO/mGC
508cwMCS5CLfM0qFvytoXK87zyHo8buzSO62M3QoOZ96uQ05aKRNIg3lCVjQkBUbIqf2OzaTrj+k
Z0Ntl5SBegCzNkPCEnA3ojA7kp/+wHCrU+JOrU6Gh9octlCZorBSbmBdFEQdpJ19KNt/AA7mIibr
C/Btia2rfIbX7rqYXuk7Pq7PtI7l586GnQDguaW2OSgIdKR5nHEPTRPh16Wpdt5Rr7mEu0IFwCZG
b77+7PYNEIPP/14M3iD0/3Ul4HLBSZF9aV34omb3uErqjuE/+xUnnNGfn6OqBPiV07PD+rtE/ved
vhGLZEkyhE3l9fBKxRLDctxy9hmB4sr/OnJTIo1KtNROAVW8GI1IUfISEXFOJG9QTtqfq+CaFGzP
8j+HtVeJ3INIlIPEQYG/yKLSkpscpyLEwQRiUZikpY6cI7qYHQUq/hbwWtzeg19eTTupXSq4xjPj
jc1NxKLcJuS81Qr7bTFsaap5u1GtQ2+lWF8RVsXIqN2enWDYW0FA0ds7Usp/hJyhILaPZIbU8Sjt
TGDkY5iiGcUmFWn2HKvQq/k2BHmKO0y+c80Z7Q9obCKdR4Fi+EwaZkzdlt7ha2Y6Vo0cOl0y3ysl
Dw8lA5b7cXOCz4ms5FoIIGbRtlbglcg9eyLQrnXi+ByKUbr8gnYCJvdKZSTjBHPXrYPZa/mVeIos
akn5Acs5rmoxhEawJjAGRhRgMmN68WefpGG0BJ2BmeBoKxTjP7uhVP6rbvdDoLJLFSlPuvUIsPM0
1mZm1PZuIzR0qqNJKCQMe8ARddQq9/Gma2BmMko8V3GygJIKt/ZzxFwNPDiW830dTQarpg6NCaHI
5NFIQhyzcxqOoxWMG0YU8RU6xo3oxnsU88AJp+T/3X7ERxlkrdD2jd6yVsgKW1V6YJUfz8Zf6Jyr
LV2qNYTLpvOqOP+QDk5/6Y+giuATsge8mBEJf5pYBYMAESLCaBtmNdRE+e3HH8KzGBUijBRnh/NO
AgseOuUeDOSiLU7ilce3mbp+uVigTbEwV7kQi7gw+APMDT1wnJV9xLHbRsQgnkYklMzH06K0hkBj
FcmTevGEwJsG4Qky0XZS1VZieNbSgpenybkixPIvWwlLy/XrR3prnhnJHuBA6ku2Vo2LAmahVVoG
UFpSG++p2/csSEf05SOzF7zWlcgjGQ5fLdgBfTJKBnqUymrAGCkJFqlR2Aedi+Y9QMWuyyXI/ePq
rNL7MSLr7gMNvncEIJ3sm3eBENvtybPexDH260yjK0pUKUJ1PO6Do5AYVAJs5h64e/lnVRi/hVMW
tWQu9T2anwYgL7EW96Z7e+PKuWtclAwVIjTZER9mhjSa8BgNNzct+igPjsctvSQXbN9SPYDqjCU4
/cubx6MjQc22twRB0RcCZBIi82HWbNfL3GOm1tjbyCP82+vDttnp17L20Epqk5MbSYInRkKTPm8F
m1RBe0/EW8v6Rfsc8/Nt5Vl9mQLM9QmnC0lDqQ7LTBq+WYJ4QH+nBSHJ4BPqNZIO0lJHGHpURmDZ
NHTrxCHnYa4vuP/DiJ7QoZEhCDzeA1l6aHxBZW3e5Vr6paUGS9UZZV7cD0L1NQykuXZViHVCwPDv
kjJ1kJ7fF/4lH7XvtYSlLCj8UZ1RLeDCpWvvLIrvY6bO1wI8tangOgnGxVAXsz4upRfvY4jbJR5a
dyDMmqIizXKVmk3W5o4eLxUWVbgSgmecbBewMrUu5jVfJvivCzL5t1H5ilL7rIoHQ5NBc6llj9hy
v83Yh2QDfeDImX1LWkiVZ98Ya5tricoeaR1vfXksMHhT7u78pfLYJB4TLuM2d2qu4tou3oJgGJGF
0IwEBHH5J3mAmeEcPD2Znse3ofwrfdTV+8YkqX3Q9unXpVaShgV0Xrf5bF1VQ6qulHvD2y3eEKua
LbGDx7I5GIeqAvKXM2Pe2ApRdLarXGk/Pam9kWdme3JoMp1HVls8rznNo+04Z8/8Js2gukeX/ZuZ
ftKVdi7ftHZZ8NpwynJ3qduIaqz7001If5uS8L1LGBJoPHRiA8WfyK4L8CUIHNVSbLubElyJYQuC
cZVU6Ka4Pwhw65j1cb2Sz1DffyU/eJ2KTEsCrkUJI6DmPcfXsD9efHWDVoErOqVwSvIkQ2NbeIYz
zl6ZdOwMn7vFPrKv1yBaizjcWZki4wabDa4VJNrgh7LzZwa693LWsbw7klqiMkK10BOueDz253ME
M9JePAk1nlevdUxmzDbxXB4XHdmiUEF8HBermE4opyraBGo3d+xaN/oP2j9tmWJ4AFM3pxoW8q4W
86Enq3ODHFC4F67tNlvwFGOQuCvzH3fFH5aETiVqnQjNKqKwVs89nh7K6svWP0Bp7afh4CruM4mA
/aYpEo/dfOImQlzdhQ+6YsVVQEMejPiwhkf3J9g9CjcJ6Qcx1oYIkcUtdBcab0RwG4+rOXTXbiKX
qfACi0dMJP+IHRVCNbgDefDUhu3g7xSp422OZoSd7JhU1bTzxMXiJvbSJkzJkBjez/qXnHJWCTkV
BI9Hy5WNIllQb7alk6WzYivS3kbKxYy/9De+30L/otJZjHm3uWjVGfzQB1i6vcJCTQwvEvDk+2nu
Q+dNsktp+d4mf9AqqH9HsjVqQ9ZEMp+0qOLbAmJufAFEmZQokVS6K+YeDt3tQuUbnuv2DsI0Rzwr
zI1oDh4rp+ThIDwpT+fw5WGyUSt9fh8xTRtuq9rFx+ZOqZA3UbphW9G1J9oCWY5kgZdm+ZfF/iql
u4B3rHVUrlEc7ULaz60RTiupobK4quz8dSl8XkmEx0vthhNUNsm9/A0bg+w482fCg0+XX1KaiTJX
MgZP2PHBCA8c3juhAiTZDacPY5tzjDpL8UW0TedFB2c8BDYTa1+7tWxYH3Odpe8b048J2y4kesT1
p8jVyTYnVITI5eWinajL+9jB2oRHJGBkQH7B/1y4f2TF6EPBjtEXCRdvnbSUE1SEcxzK3TEufI9J
3rN482Y5+vj5gFIzRL6hbFgRaHfTYeYHfDf8ndnlAKypPD9WQqjpaEPsQWIpZ32yji8h7NBMP8Y8
sWpK/6MXonb3/5dXvWnRsS968p9vmBi9xvuQlU3pAMdCPwbco/Y5jaZWFza25gdoFaXakdYB4w/h
mHQoecHqeTMC8+rhCZzLXpM+h3IQS49ChU2QUXc52/5wrTNkzV1EaSyREN4Nh9giFR94ONsSo2EN
ibKD+uf+oaXK/6j0ivzMOs5Vn05BwpYMeZhom9hwLarJa9pXiAVrerfcI8LT2sy0LXFhrRp/8GhG
t/FL5yas8fc1g5N+7uqvo5y8LkafiH03pLbhxa6rXe2SBhQe3Du8dDhYymCHMyPboFnAC4K5Y7Wx
w/zORTywKGQYYllLZIQJAhbwHLbJgdkqHr05IXhLT35OytnCqnkTNJ2QnZERgZhsFPma/UaJRrAn
dX/8hlagbUgh4KdKDj6B+SI87qZRASXQIaGAC8S1CzLNHRbOwdYJfsq4V4Yyyuq9ej7viLT1Vtum
WTy47Wf8zd7SRvEdoitn4LKXOUeBfEhMZgwQCPAFbK2C+5JNYbd7MNgOkwNpdqnSjBzZnGTVnRZ2
wVtMgfbee5m36L+7N11orDS0p7V9V9z/YOVo+5E5SchkbAY0Qu8YDNmv7aqfZEgdpP2H9SxyKGUC
sHLPgA1DvBYZCq48rV7/TSeweQBoEYa6tDx2MGrm8e+P8kfYJTdAxxkPgUhb6NjyoCFOauwWenhq
+TlykY1QSTfA+9NQsrMzBC/izQ8eDOb6wgO5vOSWrIzd3XyXTyGJXSsVbPBPliGzugPqFpAZM4zd
aqIb8L68GVnvM5oxGfpgy/HmotAx6tqLcLrVb5ocsFPeLl20bKRNL1wtPAd6xSp1lZdpSI4EofPA
9lwRxqTN+Vi1shWKN8M9EfiHJhkmkr33zDnJVbTMKN3bvuYXlsvvVK+RKWGAWoA9xhhJIrXrglsr
IstBm0VvXecE4HcnCQ/PoEddXkVbmr1wIEwyyGfPwfKzbZgCtDc0A5bSC3nof+AngghmJNsGSv7W
ln02g8s0NpwA7FokxVnVt/PgNzGJiAm3fwf4TWPRBOCCUK56UiJ518Gv/qKjHXjJF35K5i70gbam
D2kea+F8JBCm+INY2EtVf7egzicCejWFaI8MJFBUndUk+c2JIuCQhnnIdF4Ib6ZMM5jTey6xqXiT
caqGCYdCjYN5QOCCHFfiHrbXBtBBSkK5ov6DN40SEY7NykT6YXogTZmyZj9v1AK1jOu8kwYL0tzp
xzPeqpmiP/V7WIV8KpVBVaeYFjEcxA0oals95n2x+bPr3v9P4Z0hYx79l99DOThXAQ480K/15KDY
MFooWDazs+o3GIriODQ3qNuQYyMRec0gQChI7Phiak2HAidvIXoz2pd1HmiulC+AN5I557/xjLTa
gCjrchsm24I/9VR1arDIP1LybcxQcDnXjqNyHzDGmKhXXHWYalqFO5d7Z0thM7pehBiYmTHpWmtP
J1hgQ70jfSxcHuCWJbIWNAXDyzdvbE7l+uBiSpWy2YzDhQ3sGt8ntn+A+wqy7t9jjtnoJloTY/gU
zc+24nZfEvvu9pkRQFuDjmX5IoDA2+Y7vhzG2O7T6Ezq65gJyk4JLSSDiQqn6bq5CtOGFNuNSYw0
xzvE+xGkIClQrzKFiwIB0wSash8xPMUvVJLr+6uP2QGuUjVD/a/+OVJZSvPyr1a4F3HmrOmtdAtI
1DpQLgftW7eoKEMcK9flAaBGE4eZBFGViBV0RuP3SDyv5SfO1hSkO4vxMzSxYA4mlX196rtnWzIG
xKJv/wyKh/nDj5OcyXUrb6l/8ATQdc5MWlf7IQCim9mtwoApTOVk9NXhJK0Ed+Sn4GRnjO4MzzXR
zD/2vY1U30yN5P70+ssuN+ZG7guQDsVInY38KuMCiM6h2AT3baL6nj15ul8IZr/xzz0gphoZyuS3
1yQBsFYxAB3wDwuqXaO0y7GldSMarm7CdXhox4EJlkjAAeRoPQ7ppVk4IQT8iX9wLiGtfftMgVi5
+lyveP1jU2loHoaw3jOX63az5nTI7xVZijw6URUExmu9sEpyOqECPCSQSFtgECa1TMLBtOIrM7Yx
9fYylyaqRhlSAu2FINC4ZLk6Qp9GnJrFu3xG166zjH6ReJqADz73ZjLKJh1pd/fxmqBkQXfiOz5x
hcLJj0MvCppsVYXVZQd5hbeBsgdErJdKG53EnRbauI5nhkTrbNJAxTFt6BHF2DHRJuC5FwphYsTG
Gw/st5XQ0iVDo99zNH7oPex2l/mWMgdeww8QsJxAalLVpT6xfsgxM1tjQXd/s2pWZpX0ASjMowlO
C/74WDjsxtgxm6d3RUxM6/xHC6Yss3oup3Bpgf7OOoc8gVPiC+CLXv6+XFdsiIQTCW+rD4PHsV7K
l44GCpkezktMXtzhMor1tTT3AprYg7pY+lU1+ssHkW3RzPCjFMN/tExjXSwX+MejrNkzB2F+p5MJ
QFyJP4kx6Y8Jj6zjjS7uYcf+vHYcQm6NYxw2bpgNx7BzRFtmMGYql7IQbWeSKwWWGp/Qr59BI821
zGvOwWswSXH7LO9YZ+KGYPzFycGscN2i3xw4TSMjA5bMNfAGkqUmwd3sZV7D1L511YKWFE3UJjPI
g39DNTDSuMpv4vD9GT2nDOAMj8C73fAiVfmSfQOGgxB1Fm6tp7g2cWMNwcQiwQkLmduA/Vc61S1c
AbShuYrmNSTcdwx8rGijekjlwWjs1VYFvHqL0kl64fs/nrnH0NqEBMH0eHeBES4cKrGnIyy2/aNw
OeRMo4fQb9OeQAmF/ZvSWEMa4wipLBXjUCjjHaN6y0tke2Np9yYg1Jz0z+aMPKxmLLMQDKi8l8G9
2e3jmVo9CrQui1/09fwjxM29uQ4/80H8kDHqpP3emBx79laN8Yn/qfML40dtKPeSJ/F5FdEKvtsd
mwhjzehcUnPbSVrubMdMXoyC/vqDNfbkjvMx8H1NOBTCTn95AMw6X6v3NW1H+XuadGT5QM9aBsh2
NGn8dAqLA85JAkVFi0S46RdWFFOmNR0qsR7JqUZ+XgIPIfTORKOS4wzpyoGErRQ7Hokv/sBKW2C2
mHYZZzF8i4jqelZow0snCjFm5iYoreNEw97jZXfklrsDUku28D1dWpK6M57HNeSQik35224p8TfA
GbNiGb4VXwD4Bk9wm5V8IDuRc72fxpJaXqZJlQC7wxRzvWt18Br+c9cdSCnpokT4+4e7VS+YA2BN
e6EC8BnDhMuciuQ4aFpWl8qFVHf1c0vEoZwC5kVGpmWsNmvuGXUq8rB6MhkdWXASMG70TVkf7gw8
aY9Rets+Wvb28DnoIlUqaWihqMOs0kfjrgKztSuX9XnqJB0e9UVEwN+znSpV5qmaWA1Fpwjx891j
+R8STsFsSxslSIcUsqea4PsbKuVY1DIjsMFDcWdWMVVs9eZM/uRfBnFlABVcNjzVvnrYHiu96ual
F5Bzx5oM3v9e6ifez+Vbz1O0FfYfbRkAOiaMyPS9t3G4I9pxbNoOIoYTPoFBXLf8MLpVLEyYwwKo
OLtGxX7CllmeaSol2uOPNnp9ciXDcztKyrr+bExB89fUfSgKUEaAPPKXw6+xW0jtc2alKw+fsE0S
zgNL/6m6WeuZGW74R+l3VZBpGEageUK8fUisugTq/rj7iccU+mvLZ+w3fhgj1EfQEVWgK5ZR/wJp
k5Ny3JA8o3az7gKJUKnxkZArDmx14fxPL3BWoICX4jfsmullrkkOzLBLc/Bdsx4ERaH5h5nxSGYS
q/PYRk8MuvY83VB55CYzBo6GyrnWA5TL/LOTipHTL1w4vN00urruour7VGsSw9LYyY67W3OovnOr
eJ/JaQ3hlhUWzAQFRuoJ75seZGSPw1tOlBUfGdB8pGsNPOepG3yjpKv4JfvBYvQ3z6/GHPyof6bK
yEMII5CubMyFLROBVRSIq2f+mNwRbMihooc1YUtGon8JlAVMwO5+f6Uwqp7DtXAgLCrhODe4ofLm
4LYNbmnUbiFsIUqJgrKt/F/ADRBm8ChFJ5YWTzTcyr2WB0wNkPn6q7YhiJQI6iXc2dD2JApxpc4C
a9Iv1P1c+NBFsClilPybrEF9d391IMxMChRF/mJkv2gSPRbjemg3kO3kEBepBm0x8Si0ezXFKLhX
BU69/p5Am8RgbpuSCIZDoYoFinsRT3o/yLpe7JDl76sXHv7mbKXytuR5iA2DyppUapQekxvkUgtY
CaGOKDrH1gFzSNTj6YOYBAWCeGizwPYv22NkgOgDKWCF84iqXvt+2PQI29Pb0jjTBS7XL9miKvNw
iKdf5KlOEcAuEiaVS1it8ryD96FONwCUBjUV1HHfRCLJiYBxESJ0XLYcmI1J91i54d0hG5kmbvm7
VzkmgAmfNwvHrBHdIht+jMzzgXfDy9Fnmi840CCvdc/Hh4vVnWebkh4ha+nXOicjHG1aVn+zM/71
LbAChyxnKrDbyOeQ4J56WfN7nstMUc03N4k9d+hTFsfO6hrAaf142tbyoL1pTVrt6KNAfcHqC9pm
xNEfi4IFeYgSPtRYOqpqU6dD2nlmRzjrBFCIvbdDQufOcXjRf9eYeurMCqUD2zdmlA/rq7kqgGSC
ojnYiVgq9AVmk7Mm5w0zT9KPUQKF2rLhbVWFp6+u0nBz1oCCQHOAeIWOPKHz+hBW6+ppKpFU0lei
ha5gU0qHsijxUKaAk29DSe5aYwzdQhXrYMa2zTsi//hvbwFPjFk7Z5rTzkjFbqNgQQ+oRBZ87/Uc
wD3Bfh2TSxXKGtASgKXtzVQ4DMMrZ1LO/vCE+tZcYNRU9m78hJhEe0XUtIIBstL2l/IC2Ch8+9c6
3y3Z+GGaE1yruiN7VxQXsKKkQAD8SXP8zrl3sLh2/bax5gbQHcgQQ07srwXImrJJ38A5RwJEiVvk
9bt+o5/pwHccRX1NEtD4/wVWI+1+Wf5lK4OW9I4oViLXg/N7x7/rkycNewLAl9lnx16+x07PO+d5
iHB1PQopF+/QYsEpenhlXzq0FEzeknMP7uYL1rVsJdFflXSHshLZyfk7gKPnGaUQlTpe5D/z0Fvj
FCEErsgJUQYCCM+eBHmkyctNKwcSenLrq04JBJsVO+lzPpodiVHki8TuX5n/aIM/boydV+imhBY1
2kzdXbOswmKItRsp885q1CixKLoSdtLMXbYJ9CinSY9LGG/XyZ7dBf/+kDWSOSL2HkUqzr3c6XVf
K88u6EdqxKrYYgaxYvbzHUuu2n5b5W4SnAEzRMTvAXAKBGpz7Wky9odGh4XYOnWOM5ze1X+5uNaQ
KHmGAd6QaeR8WCffYP8H8Ba9ErDQ0gRL4kblNMb4nj5bvhqHjOfYGhxsBH1vImcc7Oe1u1nsmoR7
8ObMiTcn4LSTvDcbvTho9hdpSikK/e+HeeBWEhfllUM0eKAHO/MyRM08yfxjrIAftplls8pQPcKa
jqMXUsfZXkr7ZpIvlLGeXsdZybwWWvxSNk5iJUSYev7/+Vpsw0+aw/KOyv7bfl9Ebiq/4K2rylW7
ZMBmC8tZPfNck5koc9Wc5V/an2HQN9303e2sQW0QNyWgvlM4auBnG7NJDqjXWGQ9Ck3EgwEe/n6+
YXn11nlgaKoBwI7t3nkJy5xDAtThVjFVXPGV7NVi+UBOTgycHeoRicpVMWWW0UPpzW5OsZ8RHD5c
x5thOaUZSJP26YXac52GiLO+giqXXsxgjejBKYtLe6jhkx+J0pNW6Bj84Y8Eo4yKolvC1V2tZOLH
f6dJrZot6Z/Y5yzJEVXS1SPnOoF8DByKsTyvB6DP8KGYLpJOZPvOQtk7fFjIFR8GBbKzyBcXSjbF
v3i8H8htVPzeVEOxcrVQ8VvgZmE2wd8nKIjYfJQvlF+wlDAMM5L8rhczPzL0YoLGhlQG6P64nMzl
Y6Lnc440vRuBXBA5vlj0mPvTu1f9SAoRPNM5AKjZ4VZa0Sm/dtoDLlAdAUXac4ZVtmp7KLfCGCQ1
gRC8xNYTaRhN4O1rsPl5GCAcDdIrpblCImYif0mxxPFSoGwjy/pqCfz9My7P2HO4//9kwX3XNXPC
cu76aQbSNSTlKoYWRbMoCOX9+R9qd2+rJr4FB8bR3Qnh05TZvjWxCu8SX2fW+Y9OdDkzpU+BhB6x
lzH/HrGefvENwWCG6Uw6IaXruuD4MJBCDn/hiaPKPeenZUYcuESmTVYKSz4F9k2+KMAVwrQFGMg7
C9vkyanxUuq1AFlKlhS1TLXB2wMAOCRxsUq8CtJtEs6ChiUQsAQc07WSn9Lm7Rs6wcsiCGmhYJwW
ICprhytX7lbYUoW/hrSNyqVsZhp+fjLvJPfwavRxJVLkpbOwhjYJ6Ob1WV6b8YzLMhPQ57SQDs6+
/uspJjL3aR5X8Nu2theHGDfu7NocRpHMYjPgmzlVuayxiVDxLiXEDFSYe5E8Yl+0q9ZlrRENBuZL
2um1wEf3BWIZwLW7Pu/J1QywyHrUsXLNLUs3zjaMv34s85670uFxshvR0tWmYTMox1BxUHH80cXs
loAZikerlVr4J19CzXfzVbo8IQhpd1ZFKRidR2NxhaTBrSHIyG+rgSJ64YtJhkl0bmaz21Pdf2a3
5wBrtQ0Mq5q/MBtNSZ/cH1kop4piYjZiUzZUqP8VhlAsfBtUQKoFPmwW1TsmugL/foiDm+bVWkC4
IskgF2c91gjOSSqvjRNCnP5PKRerCT+FT02FfUdna0jjtn7KQT6hHLhSwBL70K8JI64qYWgWyGPO
t69d/rKQ+9kdzYbhGE/FV7q6xzPp19T+3B/TtnElslrJxBKOURtdqJnPJKTNY8CQBs7SQZqUt0Hv
/mujxq0dQk5VGmHiw2Xxd2Tr2yto0aCP38lwuUjtEeeasGBtxZtxDQ4+f/DYAm3bWumByxSjddwZ
0VozeSDv1jIAoo9993gjAgqw/w7ASkNTMm02dxrjXXBqG98EgcE+tye+cu0louX4QsvUkIzxTWM8
TTs3KPVkWK2oKX69TpNFJVz2bb6kar1WQMSaObUD6bjaiU8CTo3pzkM8saO89Kyi5lWyinIqGwMB
d7KIlV1ZZUw9wIKR2h0eNEl3ERBUE7hM0NGChsykEJoz0c+6hvJDC3IZ625S/jTbb10YGI9pL91U
iRhrOk4mwpwEhCl3la6aM4BsX6sveCRvKbVluGG10YsZb9Nu5B2DAE71F/pk/EvBUAi1Pdi2elJZ
FzEVFk6t1gpQQZtrQNUovGx6pMvQE1w5rveRzc5mr+CPS8Xb4WS1fLPHYRvkeaKy5EoxPjqWnY1r
PGObMRjsP/hZl9iK0IjPaxOprjmI6Q7OE4bKlT0F7xC8raBozgIt72vfM6dbw1VveditYSlERJvO
3pV7/998ZIfGmYmAenIQBJekjHGagAm4ax1Ho8BxJRsd+uop9nz5RBN1Lbi4yFfP9yCSCRoMw96x
5z7RzkCG8luGMNhwD9hwQx3l8Y3Wk52Tk8/d5tkrhzIGo6M5uFdAWuWusG/Kvd8tA8nzhaMmYng8
8mgleREnwuFWvHg3GO/x7bKG7IYw8CYDtRGHJXcwAqixuEYL1cO/MGuo0hzAPcv3vHL10BXj8DyG
dTEMMSUWygxZQu7n+tOzPmsmzS2DGgzU9K+0PHAeN34Wqeuu56XJlL+MxcIwGkyj0XJ/PWiLDEMC
jyY4SbHQFAsyGoa+w/bnzh3SIMShdnYZYG7Fg7eKay7EKAsNqo/I3r70Xd2MTjN5tSZXw4h5bqW+
wMpiAnqWM5WEHC2S05MNCIkN9izj7A4oHOZfE+px8rGS1L56Y5ixWVGtnFMt/wmO12TFXheUHr0V
sTjU/4rkZsi9Lm0gxgRjUQMfrgNofWrUzFJ63unBYAk9mHjAS6Ob8Kla8IBDJCYdPquzjdbmo6fQ
Lof7oHzY/LTFaWbAgI6vXcZ8QrPikeGsVeJeyWe3PBO8ZbEM5RobzjpG3tXgysWWIPm79uvUgobV
O1THXkcWc9DQ46AucpAauLIYkZfk4+ewhv+gmeIRD0stL4dIqNGlva8kT1lK6usZpRGPNIOGnTgY
8aSt5NoVitMJ3GTSHLGB8Aldku8DOtE9xYY3pwwQcpEzy56HDZT98ho7jTvzEB3AN3ozu44nSg0E
M6rv7CPVptMElw92RifCj9WGjcyLQmN/Lz5yg9ZdsoA7bz0jmPVKEm62DlyNKt6PfLtir/mQ15su
FXP8ddfmysipWRpgoeZehtSJrRYH0CYkn0zkgF46KY7ElqrT9nXB3af8w90qgApHmzYxA10kx5CJ
4TjvHwqKUtK8oABvWslRg5ZA9Nr7LxK0D7o5OLsenmd9nTXKZtOXNKPrzu4ftkPJ1jArZF2zOSJ4
N4s4LwJFLOGblnhGd+jm8S6lQSiUxA3EdKZQw5yuxfv9hjcTT1Y1TBOfP4r2wiFP5TBBTPBBX9hj
FpdELhClaTHOAKq42ko9+rFLaBF1mINyL+dxKbeWHBMVX2DhVpQHGmsMzMvL5v3IJ31txt7Mw99z
jB2TVtusF2Y9VgelEVVUKBw0+OjDMHyrL3YLV23YuxSm2LHOxl7MD2RVn1Iu9NO2MlO7RKc28IBX
Q0pPeyEayMADS3UykvhtxkilTZxK2yaB5yh5o1l1vBwah+BeuxzL4ML/j/AA7Eai4k91I9gA7Vj4
VQDNUvbYnvNuCxkx3Y+HyaMYIkO0GErSxsTf9yFBqF8nxvCR+rTaamPvCy/WxjFvtFgR5G8FfKNO
ppr7CU53l/x5ed6CEVpUW9GQsQvGF6Vz/yg0hluqlzHrA4ZCbvXX5sYzH9drh/fgFw9k11dzTw4s
G5sLNhr/8/k+wPvwy8VnQdnqEh6KI0dwfO8aqD2WM2cdk7H15+NBWBzsmk41wALwPwyUrTPPmZAR
T6tDJIlqXRnz7S+ky3JvvfAjEUDboRlu0nB9IUJobeLKwenynS/8gBu5Vgg3+KdPI3TAcFJVadwS
Pvp62kp7/Nvhoa6u4gYb32PtmT5QHH2LZzul2j9Vcf5wQSdnP2wdZw3dPjBppfkbJbgD03loMLtC
iOcbk25KzGvbRogUP/g6vrUSh2BhHQX4LEcwK68SZ7v3xK5816VpDGP6dpDMg8Dj+KZadep32JEG
IixAC0146KO5M9y3KCCczzrG83rRfJS9TMn3G6Tfy3GUm6okG3InkYHrXe6AhS1r+P0QUUXYr9yy
y+ImzLNtsOqYJL9WUE0jeLcRty9EbJ84kSxe0RDeIxc7c3LPiJPNjW+9OFqOsQCP9BVw/+zqr+PK
QXaHFXQ+pNlD/aHjL8HaEghO85ulzMc5q0D5g3ubdG1u/bwH+Y4s98OIAznDnL/pWkZRkb9JoIca
HB9k7GL1YnmFWNAV5O8DD+0xDNZ75679y8eD52U4LZz6ksW848ipNHUvn6yWRLNwZweNSy8UC6ZK
ae4+9snojX15v8ELMLo9kqKWWv56fCoS5J0C+ToP+9fI8RYpP7kOtp7nNmY9mJfgIsPeimCbWEHB
0vz/w0ImmaI5xlVwDuDr/e/aqZKxCyP6NVNkkA0tIqnQu1jHBOXIoVyTOcYMrWpKHaCHP0Mj37TL
0DSOFPffXiKHAc/MbxPt9KrzgQ9E1vZln/la6TzXo6ViDR9RZRyNZM+MIlKOH/hP3F6THpXeztX9
Z5lHRJ4BF6Aff2f6UQkh9d/aSIqKHh1vENer9q+jtSV84bS4mVTDyysB50l7eA0jeFVFWNBNzSIC
eq18W/wd7ecfCKnnhvkX+AQp6P0XjUhohTqL0Z63swyKt5OTTl1frmiX+M+FAcQL6jAn8rYF7c5p
e9sq6EPrHPwOor/xmKNFYZo00rqUKAoHUwHusy6VFgH3in62cAVZmyU4/1z4M7qIH/1GOxrxWbxL
+C5mQxjPCGwEG9IKbNlcacNhYNHbhkUQ6sz2xs6jAWsCtequHqOWGW/6pfGOxo3aKlHcPIEcYDlI
lR6KFW8arFwl4lFflPcF+mqHpxl1UwKGoPGUXQKdnxNUAFc/8qyKXSNKBIprwZ32RB3fXXXg4u2N
VtatEokokLo/f0lNM2DzQyDEnKpqwLEWz4I+owZQunFnW1b4IW9KK6I7yA2atnnNLxhLRCg62TDU
lkfsGEs3Csw2ACvyzM3tMWcsTMOTl8Y1FMvWHKwuL1uSS9XoFI+t0VkN7BRHYA8qMnaiUAtYBeFK
wAp4O/CMhVhYa/98c/neM9HLjBGuaCTQPWJvpvpszD56jNjNAhdjXwCRqM42UR1ILw1IHQrBTC+j
SZjo6Cig+IXuHAEdhJF2ORb0VTur2o+dVnoU88GerRersv7Q7QFvkVVh4RqhT7Ual1ZWSrSwn8yT
hL2eDVdkITC/tf3yBrICS2il2dkK8vFDcChmZCcMy58GqfKaLB913DKbcTgyskhFgFYmdhibCrKJ
YmTcANlO2zA02DHWyZtbGKgtR8N6jMlQNUddUEAGeK0B1yG4Pk40BypJZn+1dZ0boMNVpXJ6q4cx
Tve2YsJwtrEW3ZaL5KyP2vI98ewXDZs8P76B2KIbqPMVe4bMShRcM3S6qtfNzVcnDVL1DgCa/xWB
ilFf5rt75xTSa79xsE8Qr3IRw+kUQa0D9FFGclfjEGz1mnMozYs18+Tgg/TUO2uAsdG/e6t3Qogp
fok2j+H2iSIPEvz5CrCbszZyoOORCqyOn8tFR6qhud1eqx4pELAqLKxB3uQQr8xRGiU8XzWfyrIo
xkbd6A42Ep2pAbGAJGQvdYn81NdN+Prli6bGVJ2tSEeodWgyhsL4a0ZY8y+8gkmkL8cV1g83xJX2
afsP+NgE/qs1g08j9bVYPb73Xl2uhUzDkUhDXj1o///NAxDCjsOZFj2B7aYbprjHutJIHr3avNKw
Kd3wJytaZRkd231N6dsHVV0xO1G8DuId6tQViI2MjHM/hOU0xr3putyZCun88pLs42oIrjbBHq9K
SyTGMg6teprTe3qD1c1UtCKM6UcOUFJ/ERo8+vot7Hx3F9PblWzTeVs2x5v8tzLuv7FeHOtoR+R/
gE7F0c98oLKKLoVqIyTgK6Ju0h89RdlzA9V0e30v2cQp7rC+NHjaoqRbDVevexzCFzf8p3Wxn7Mx
3QoEwPq/bnjl9Ve1aGxELKlRgnI4YEbJLdrBvfkCZBKuxnvKw1brLfiaZGjqLVvApAP23457ImCL
2Tq21ic6J+xBpfLOMlxf2opmalGuFpuzpc+SFaG1qDs+CgLFnmokh/EyvdJBnkW2lkncV0eWOwUz
MNrHGeQ0FToDS6m96BdtT9Rx4f0oskZxpaIwY6100ceydVXqwUKqsnzL/yyoQye8sIHAZvcZGmXM
OzymGGMXmY4uKhhP8jOGej0DPhzHGXAtx5cOysS0xFHlMKfm8ajK0lOUNPsF8FfU/6f3nziJ75AB
eSoN+tvSD+Hef5lu7O+T8EdTWRGhLoezmMN1MCeGLCeVaKOOs5GFrqykLTtUQQgBykYiassXIxLG
2iM9QjDgjXDHX/jmXi1UETEvjiocpMeApKrOVsreXizlyThNtI0Wdhvn+EiQ/Lagj4kCN8rVoq7X
j8I7x3nx3c68RgFVOpZFczH2dpSOwd9PMYe6EcLDL1kvVE1YYwSx62ZOHCKcu8SZc85ZwrCUXxpm
c/vwgs7ThySuiQsx+6NAsaQLwVxZTNDU88WcQklwBKsY2MnONQLEvLekyN1XGn77jfNwMOiKYBvA
R1no0s+6JWAunhEZwTkxl7CTIkdE3YOo3J9K5xMkxFW5BqfrD2AfNTvZ/uDq8QbzUtYxht+ZApMg
6avtUlQpE0ErfwrNWBvpZ8bx9d/vf4dMV2Ah8nItIW1Opwf+nBToO6pyKl3+UfL+em9nl8eqPGKO
54DI2ZhCHX1vZKI08cC/jdIM2YUs+0JFj7nK7zBF16x8O4+ep8OqXnU7SNFzXCL+heRuaEJlzE6N
zX6pTY5h/aRteu/peOnc2VksvxjvWh4QOrD+q8HawnN8p3VTr/zpWPGAsqQY2LklO1Afm7AmKOWQ
tOluYnvRH9U1k2azzJynfzgozCEUZjz+ctLk4lX/bCmAFbKP6AnTyg9ODVuwQs/5zHch6Nr+IglV
7KkqGXEPTt3g3qMnWD+JvOOokV9VFt6UA96ORjQXlO02QaUfI/rsc9ZZ8r7WTWdFAztZZgMECKIr
cS1LVgq2vbMLImN8MFEKj7yMgr6f/zNO8YPdK3XIuocEVnJaW7YNztrpCUfkIn9gBr8tFxIB9b8n
YDCiTOft1bzxKVIaw7lsINBC1LBn+YtOG4A8C0bRYiF386ZPrXtB9p04z7xxO+pqSY6T9Iu88w+i
aGCv/+23TmgXNqUJceGhcTWAZru/RqygW/ER/mQgIY11H2RNwO20BU1xYN3jeQReFGUfeL1jBBce
YZs0Yjjt/r5ZtxdfH1464a16+600F9KX1o0LGscuVMPJJ4v0VS8EAas8CIrQRUVKW3Ty/CD5F/HU
J5NXEsNv2xpaLTPTwWdk7Ijx6MkH+mtCLv0edrckgV1h81PhIxsPW1ckjpbLZoAz2GuubZIANX9+
XcVvxkYZMWtpb85HuwZcWFBXBKenunF53+GaY5F5QzxFKREeRBoP8pm0h8Jym12qQg1n8a7PuYHt
jw3eO5CsJdli9zDEoaq6GvX9lCNqaCedMxvGrPUVKCbGbxFeeif/83yhP5UFFWLOj9riqEPBKIXl
lm8ZqyRYfslxn6Gd2aubWQRbRW2papm2Lc9E7fDys1w4szXn5JGGeo0R3IfbIZNGmSDrnBJ/gTYv
6inFRj9rF8mU/5CKYxLeFqyzqvnnvMv529nRQOSulWO3iq+glEQMaCWloUPJcQXPetiDRbiTty1q
bM7K5GY0G3/4AD7ABEkU+AYSj4DZ7QCwhKxcW7/dsgxCIrvbX8Rw4OpiujGhR51fAxc+d9Lmk74g
BU4XGEPUSd2SzjZKRH87OUpeMBW1qVcDVRs8Vh6P7VAlDDLwCITQ0DjeGZ2HEjPB9uRjQRnfgGsC
6Y/PW3D1oQO8roV8IDxuyS0IUA7k+wEVzmzD77pBLMKhmSJBJWtXeRF8eH0lDsuyyEqdo6+0hvov
U3+nFa1nGQ0v1blWnwKQRmv7cH7JcqL6aIYUPU3Mhj4eEO2uHKCSwz0AB/r5FWjxZd5kpdQoagwE
Fh6uZOt6wWdIjp2iAjVo2W/3tEnMctRWCEnn+dDZbCbuIdwt1QtfHKD8eXAucZQqqsKXyv8ElNDq
Dk3NLZVsDkZYsE6qMhlg/cyBciLRfmbekjrDD/F6CKj+D/Tj90D6AUYK4Hk/NqXkQLTT6qBQDfKX
bfOj5P6UCYfV4GTejdeWbEcWExJ9CS7dI0hGuaQ/xWOc9Q4eqX6++xLqNMcUj61LYWyAjlEVDxFR
R8Cjqo9mlbqMSoFVU5GmloH04GeylIZmVaTnPLrldUm7fa7cwey+HGLwyEWFS+gdtHxgr6Vx1et6
JfM+GI9mGgQDROw/HRqrVVlxFroH4beAvqs8H+O3WiMNYY0/QBpac6lgmQtidoTsm659OFZMLuDa
pQkrEmRbTibgPtmKRQcptO1p6aUBw8pPNbnQJysZWa1kiI7XgZ0JcRXu0XQ4UtY5Dr0jcH4wKRZa
0w+M91Ye5uM7NTBdH9v9YvmWCvtKwE52Dk2rYyIVQh0YIYEGlBZX0OsbC4lVaR4kL/AeZwLDPgLQ
L98KbeHTbZc/fq8AhlQu2k+cg0h25qLASS8MRe0E//feG4oFjhTs3aJgh3yWQNbXxYN5uUas4Znk
eTx3ciExPf45VJIAFO0H72QW+o2fAlXp1ronvXSoDuKupRZ5im6P4DWSHpeNCKjW9xRfM4+WmpWE
eO+culM7dMbimIV/yzThwbPJz+ggcwUbx/gB6jupon8CzncZzomCh/6grOpwbHuHEsgCclQeKHFB
88slOxvHAHPDsr5SdgI0lwaUbtYcskdeQ+CYLrtchaiJLuyHMhCw8iv4QN25BSkWP6yywtfjeWxx
d8HQjkpJKrwrxF0oySt6HecgSrot8cvc7DQP3gGr0rPqzkZcs8YPlnmHhHJq4ly7WubhFqRTmOv+
WvvJKUGGyhmVnd+E95x0id0aryGBlJnSpFF7p7qkyMVyz7QICG4En4frK8XzAw1OrdQmULb9cU/X
xq2S6Xsu0xkYZt8IBQBZXLGGaN3LKpTwqKZie8ChG0WjVWcJnU2jT6TayJifjE4FRgrdJmsH2Ttt
mFdwhjAA1YURNkM72nLeW/p7Ih8bxgaEpKQ/aLkh6T1LOOxnlX1f92PcC6ZZs7UqqlBuUsygQMqE
By1lhqF5MUNpR7Byhg1RsukeZMhAGYlWDn4AJWGvoeZCxE2YvnlA5t4lzGHcbiuMff9Pp+5nPxUg
o4KiSvjgTd3xNak8uvkX6fylIU07SuvQAOf+rwQx500Vl5j/I4ka2HIr9V2HshebPP7Ns0ScVXND
5HPh1oqC2cjMscpqLDAdhDWN6Dvn8u3ZvQEaf5Ijxvkui9h1Xa5/7Bo/LxMEjy2Ojhoip48K1bs9
Yp6I5mhg5tT8w24w0E5MVaFwib0QPFD+/+FD2RZ1QqnmbyJZgVO5Q8SpRgUu5fbp73zgSFdhQo50
L4h5fuubJs32pN3RwrxngRnFv6Jkb2eLDIrd6zmS07b/emH8gDWh/NHggQc0Q1rsukBlAKsCuHCG
o1wGrpdopsDLf5ucO9ezSLcA/Eq0s2L0dojKJYKJoVHAr3visjbFDJEsljGnP2njMyrlLlKtpkJM
OpcQf9hWBJVNOspHoGtCHEmuXCg9ocRp95Dvs5WU0M/r/YHgMktgipobh2vOUV+2ZBKy10PBU3vQ
7RAijxxtcVeBORcdi0+mCBWaeeBjDbf69v4KyhAOQqLaJ51O47dkoc3mgN9gC03TbZY7hzxUpCHJ
LDHDL7GcS3X6M/LRx9lnnCxo4UcxwAllZzPkbtZt6U9O8YjdIxZKicnlU2uPX0/+JD6+pucQ4ChV
RBs5UBsu62PpUp2VHkh9hV5xG7MAhH2MgOluHN8lEl5sqftmNWUCYvigJsbAxnPTuN+x0MIXkYCl
1U7/6ns1GwM5J84H7lJh9o08sPNW7CqmCWUbR4tPUkhFZa+ALr09Y2ewgnI73zOENUbI7j+42sTU
esxljqoF2ejep0cHH/jijUmOiNBxCJXDVnflvvQWeoywkQXqfwbuEaH+vViTfFQBsshV9ioF6alr
GFx3KZc0NUKRADVcpwUTRh0DqzNsry2CJtTkZegtM/aKdMKY2NiKEvYQ8Msh3wQ++Fi7tf4j4Uq4
TNuTVwzPRS3z/TOK81kXDb97mdk6u3/l5X5pQttz1L0DV2kGNLDWTN7ZrhIMGBLzdk25wCSh43r/
KdU9f9oCFYifG3KKRFfpHQYyeodzbn4+Eaw8Kf5lKfPCyjXx79u1i46Yysg0q0f4ierhl/hhfi/i
Hz66dcr4ppZwM/xplVp+Yh8Wnuvi7JTjZZSikcEMwT4hIq6P5Vv7541N3YXecPIQ6kUPbKynL4gD
4YT5jXp8/+T8a/VuEUuaX4UQ9foo7smLKm72TBPIbcWDRFy7G4vHc9RhZLK8f5iYy3PsrbOCiSit
LVuQ2fyHBkSMaO0nB6t2F7bUU5/H+EmTDgaquv3N1z2R5GzjKKNZaE/sn0CTnK1OR148Grf9vZKd
pdTef4K12jZkbdICddCUVhyeUxLth137HLFi8vUcPbXKix8g3Py0RoqXSoQyvADWfLdf+zHjlS5v
8iHdKJAUKWszDNjvqOlPjNzoBtMZMOaFHruxzsojySMNFiT99A6O7ynZPeRBjGeP6ZBQogebpoGC
V0ws/vfTGNejwg05RyW4iGT2FI1r5E6aiTrqEWRNO1LRTrJ7kA32Vg/slXXXLde9SdbV0yNs7OhK
twd6I8PRS5F5xgVMAFIrHEeEbd/2sx7RqQ0d06iZmD0d5YR/m9n04GUWAeihOQ0FPfegzx57E1wN
iZZFHXBK93KC4XvAW3SXfDLnMPy16yRXPQhg/5dAoeiJ6mW6spjRjKyXy8+/nG7zZMZ6fQrmxrPz
fdJV1nL+NL/nQjiYVUERbp0XFQZTR7VP8UiyCdpxyGQBFSlPGt/STKeGrX2NRx+k/YA+yrmSEY8a
7QSRuf7MLdYUdJQL8aJcn1S8X33LOuAM46B3xKgEmlmjnaihWquDykdUFq1Bzi73NTvN3TItAjxa
zyUxJSAS1rnVBsCExvKr7eN1r/n1kAsHO4D4kmr1L10O6QrnhNOGJvSQIbQjbq/dB0YG7AkI2lxx
GqY1rau9LGOiHSl/AmgS1dXHf2OcLHnpwVhmB/WwD+YT17Gp6Z78R3F6GohRhmuwxKTmuze9zq88
L0GvgPcBjxaFEVa13eEpX5/MR7xoPI8iMFt3YZ7aK89V4yfTkwzvsYXOp4vhV2cQUMBwA74x+XON
1KHuBT3EhPaNvQwGJtQZQzw4NdilBS0TDtWONSMdqYuaLb3DL8DG4csRPSUP2oJ8xVXT0v+xITM0
6EaiNRtOEz8PmYmToryDEPbaYQR+twD08CluabIQ4JZ1SfnP68tNl5KkaZwRPw8LmG3BQ1OF7Xm8
KUMuofONh/TMb5q7t4//9iwrBlY9cRrjGv61lBpHrd546qapskLlKKZ5S3cxIKmV1HR9l8hmdhxT
Obct6wY2cJmTtt1Ve3W0n02cpystnvCx+IcjeuUXq8iRDnHsOq+Fm3wpiQPZwK/DLA/3QwqW0QxU
6bw9bi9y9RXl3q5dlSJPu2XP3NeOroSlBLxQPy09hB2E5Jwb0g9jx/gfnHG819zSJ6S6m8nh2sWr
h2npsAJ4Qjr0VgV9yRFo01xbYQAafm60zWVhvwWSwsVJ6tA+ZyJWOSw2221cmtIxR2E9v+U2Ys7D
bxS+Ao2FGtCMlrRAGLkodPaYkOsVaShbBugljJkPhzrA6qudeE2Slu8/zBgQC0VzyTuzIbLZcaTd
0/QMJKB0ciXIyMgOUQzF3ETf6jDoqpdJBpxDx8ih4w8egBLhNGcvcty3GZFl18RRSPxVeW97Vdpa
d9fhzkgLMGmAmvak7MeQ1xqp2jqRK+9qpSrNMe0edgv//AFBM0Cqi4TvdnnKPxPQtwKA8Djc9KAn
OF+bbZ1Ue4NoYLziNkGc62NYBMQD7iElHztP9cuEEgG+RRl3/Dk32B1QNOU0mGD6udhcsexBT1fw
3CkIbL9DsfjudLlsgYPhQ1AE0Q4E/dYUIysJQk8tlySnYwKAxcmYKxQav+PhyZRC7E/8/TrTDdKi
IGwUhbBNEG88vJ4gPPXWcUnYauFM+2VfvriOpvA0jjux7/ijMWu4XybjuR01TATfWZIXBRz43e0e
mK+IV9n2qA7uEQGhpjtiNyorxExA8OtqSR1OQ0WZsyOecDUlRURDNHHYWOdjMvr7/X6N2nH3v/5D
frgfBBD7AOd4ms8zrkabCrLpeLPMJNLjYwl0OryTRAYnW+FqHORF+I+HcdUXybg44RKBbq3KwxCR
bM4YxKE7IaUP7dDBPHKJViPkS0kpHEwEFQtywhLoJloaNtd01iaAsRBHrNRV/9XJW98A5odIi+VJ
76akR2KQy3cC5LdanHIiga/fYrb6jxJNcQDSg5Gn1fjUPZO4tkXdB5fG10mao9EWzacvfo/8+6Xh
tukNF+EpGSu0tpZjYJgSWRhfdCRsxBmV1TRcks3oEiI3sLAuKm75tdRF3qdszwoMqAZwV02CXeti
4rRL5NmOQF9gLuZ6Hu1hZ2qbLPisqUDvWsKBZZfAuR5DyRX/E5QRRFM7/ebrVXXQ82ucQDCiFroo
nVSMfVQ0lr9u4ULI1CVpj76HBPEHH/yQwFGyxHCzH00LRQoQrHjzVX0iFCWEAZPeapqgUReWpOOt
8d2tLpa1MLjVeUi9771RzDQd2GNuNG3hJPEjk6Ov7pK9JSZ2fa+aGFLBHTr6M4MGcUy73akvQYyz
WlTvsXp7OB0fJUHLpm1bZI3H0eMXkuIV8zdKIxuzyEIARz/ffUllPGz41Yqa0U7Vd8/bjCZ+6iXD
y4VGOAp4W1aecdpwo//PyW44oPFj3ck6tQh3kCjjYEBKRy0y5TFB9WXiuWOcYx5h1jfM8FQGpG/V
NbuLmRe99oaQZtsfnB3YI/kEUKcKKttPqGkQMmiY9A1ruyEn8oSB/p8tNgdDCXNpjzwgzSapMBv5
lXaOpmDOdTV+IITvutNmU4x01va11bK6bFrxRar7Y0mu7d3zNz6RctvnLcgKJUYO3HXgSXY6G88G
XDlGLPgFTHL/aN8kqHiB4gtoCg3tVe1ta4wEqZ6V0NNrGi2YG48YzG1hjQeyJQCac1K1vcUh/qNR
K4bBC0NIJOI/4gc/dkZMfh3RzdxvIaTANNAQ7ZzA0XyaWkVXmdtiUbQMbaME2fIxhE7Z/CBEQ9gQ
i8TncjMSWTZYl73jIV7brsvXGuRexnTw/h8o+OHhotzm+GevGBzwEKGMMXE1fNNoiNAKzrZRIEaY
7kTEIcKra+MJf4tp96WV3oAbsvpcOzfZN7pP0QHe+CPNP8c24wcABm6Hy4Yac6KHSsC6l2eQqOKM
QxESNoHFg+fDbOo2Zn2H3zluI9YSXOp9ZDtgEM3Wvz/JzagOaUr+WjMMvmyVMBEe2rGHe1vgKrVx
H4fNNejHxuURl9us5DCTk5ictg6VHAZUSnCjNkqET2LZOQ/bb4gu6GObzM/weGCF8xKRyfJ/2vjI
0IwSN7/n2/mChykxfCSmNkSHPM8zg8Z8HSWeqNiZ/GLsRYAJdCb1ir1j4o3dVKTp1sz/TwXS0nUN
1bCArPYyIcXnPPpQ+ilUWQpzyETmrvyVTkz8yBvUdt+spWGcE+CFAGs5/TKvPyhJmB//mctO+fdZ
M1sD9yx9UPBFRGCO9dOUYKXqVmrc073+l3Be1F46N9T+waLtVf4JdKbMnfIyJDTLCwJW2Qw4Lg9i
a2ljfQuaMoNMVsLcBAbBxbxxuSpD8EDbmZKs/tAa1EHtELLNH3msrNz9Rst3ITveUdrcn5hMF4gU
MJZV23OGDChHrnh/6ieMUJHw8CiplR9xZRHT2rP7KwD9oPBG6h72ykomMHivf2jZILJarPUCF9qT
rZ1ztJHoRN807AoRVR5X3CxvLh4LY3/b7RnkyH8tln2J+4tlwYZbVdo89xUV7YiWoQ09EEvGmYpN
Y6eq03mlqHhQQTusGuW+eSwFEbN8tYG/FNxgxkh29amDI7mpYXWth7TwtdzdqN/hY9ifGi68AeEQ
nTfkseFrQEArWR1S2N8m7TcycKYAEb+y6bZONRGG34HYoajl/ioQgOMfuTfpb860UGfEMI9yUDh3
+FLvzNdI0wC2HHlUgm8Lc322XLJ853UfPNWVST4L6q5F6GInWnd0y5Pi4ke8yEBEOgq1GQyHqZ+L
a50QfOh2ruv9ifN3fdlEefYpyUbFLyrhu+P9WBru/TCKoL7GPBBn/Zsh9sF7+fxN5j71zSI/KALa
ICUwVB/p4/u6/zDozZIxK1VItooetWnFoNXNnE+ashiw/8+oGrgTp8Hy6/drs6ephh4NHYfDpZ/4
UdECImWEb5ceDxZE4xk06yBVuzixRTYeEBxFoFvxWjJy3DQqNF3j1zUcK2ddOvb+lavCc+A2R98y
LCBdNzfiZAR9qojssKHMlX1yWjzK7tx0cWfhob5HV1JeJyccSSEPiZf6VyZ6bK6mChP27gtAc7J2
ffro/+vR4uS7gTv3wGUOjGkP3Z2wY67xmIaiR/o+7xGKm0ObZtWPkhqDoP1tOIPaSFIMFLOmmjp8
S8apK72x9oLka2Ef9Cpao4HllzIH8SCXiE0Hr+YK0pRkxlzcOR10s9qpSF30OHt7z9kMPnpHSjMY
dEZWtj8i0ujIdeADRwETxIZlKiz2ZE6Upf3lAYSqou7Gjve0JAZ5+SWMQkVC3NoJSMp9qyAUuoul
mEkE1YkAk9nwManeqxKV4jc1k+iXTSuW9VsHMmWsuUfLy7kf9vW4aBZPsW9xuw7P+zHd0WuuP31Y
Qn6NIs17RNS+MHRodschkG/Sn9rBs4Ubii3rDwB0AOwH3uaqQ/8WYTSDrEhllFwmrDMywlxbcg/K
pX4BCiVEYH1rhoz0UKYzIicTtDJ3Pg15vZ+Vl98kd3gPlUSPfVapq1k+uIfT7HvY3EMn4BqtNc5i
VyAd03f8wdBJy9ZgtXGhbGd/arwkJXnrk/qOrkHRjAKmxZClSF2tFTDs00vW1BnUCxr7k97EApXw
e1f7PBGlCEqZ8bFAMYJVvD701ghoUo8SNPKPwHA/48fYmB2dTeGnzPBfGjLtkA9pTzIY8PHzujBD
8adtqduMLDRzDibY2y/2Kn3pd/ViVBULx7GIGyt6p2xdd9GUKNVuRgshI0VQrRK+pdmEfQysI0TS
aTNM59xMFIBkiHJF6W0XPBNvlrilfnsJN49ROCSt6W74YUDBX+TTSSTBz5M9xAOdECvbxS++QTm+
e7PxGvTBJc/kbgW45eaKePpILCQzTCsDAUWD4tifRvlYTxdqQfzeXuc2AFsTnO9PplNq6F5G2Wh5
d/B46ijo/vFxV7ERnPkqw1LZmR6+EF+DyHvoI7Br5NWIH5ZZHdWafNLtYPBOoAiSh6yPVobHpoXE
fqZRxJm5zNlM5+LI49KRBsxRAUfZZwTWaw0lbrMUqoi0j6XceViGIC2db7/PM1ZLyfXjX9+VNA4u
Ch/3fY0DPisRs4SVD83E54G6H4Te57cj+/KspvCs1bej5OOya9fAKNbqYyD4Yz7QjfYUD/qB9t7u
2YWWuR7dPC/q/IGQuerQ5BHeRFURycWeuGh3HScPPslXbF2+ZhS0mBDXdOI38pywU8pJOdz01ROo
OlN8pLL5ULN8iXQG+fcd5ISsq5HngwNTEyKwtJctsYmf5D/+qJhf70QMIjX19Ke5XiJK7HF1fzqx
CBqdq9GIJmpBVzPWLt5dHgMzJ5CwFA0PKEGB6j5hQJNfLz2Od7/MaHqCZxTVHSGAPUlGxuwB2AJa
q5tWxubJFN7W18ajC+MShSWSUnkp3UQ01PQRfzBPbljz72QfeeikSCS5c+4BEKESXyCGdkhDblWb
kvsEzSxuadoLTDqSOOzN5DdqkfhtO4gvTjERiqjmYp4SmQoZmlZ9px0OYSyE69QBso33Fr30bCxD
OHa81AT8019aBfviapjJvQTuIBWtcZzbjpsXdWcOvb433Xcq6lDyx9R1Bf8iUEInyXNQAWp4Y295
hvi7SEbWO9X7hadjMMgXe+Vtc0XmYP0OCEWO3hJ24hEWqlM0Hl6tN8mppRFgB1yALoViiWtIdV54
N/FeLSiEOWs7pvJSmG58+Bvtf+/js90mkWq6WL1VdHkdT5KWU9NWKC28EQojZpguy17LXC5C7l/2
4LTh2uh5NfCpXqTuaYGL3P+oBURGJ98dXF8/Qh0Qy5rFB6ozbpOeSLNdRTOjV433sxpJ5VIEtcnx
Y5igC4A478SUMJ+uRl8EjJ9MObQ4jF0k6jWjMf227sz/AaWYF48qmqA0HhW4UKFGD5YtomcPPrr0
kA7n/yNL30GKvJFDIz49N4SNkCzztgUE57tZpmmKTLOyggOLVNAJrZY7qpwoQMksPLhZEqVAAjuq
FO8WQrwjh5McJNz9B2dsSacMjEzX2Rf2wiNBRrt6J5WdXyOgV7JQb/SivwCxJfEbb9T7AyTkvc7w
8djfaarwxIza8khubHHxU47CBMNVePK+zR5tbC+h4Zj5WpWidZ1N90yzDAkFq3iadFwH2nePRDzm
57JEBjA80obSQH1P5GaeSCL9+VSSBs7ueuMAX7zQwo21qxXq+y9y6kCvV44tZp72ur8TyvIwX3Ax
GlJTjIISTdYKYKky0c9z1x2hDQbn/VvZXnV9Fczs2pwj/+Ik76kYoazq7Wqdfb8aUwb5meOQwNkx
NQDv97oHnhbKT5gZ8JLMcJlDxSHm59xMQOhJuyL82YGzJe318CdEZOXUV1Iu99WVuooVsnK4Mqf7
uPctWMSVuW50EPBogwZmP4hY6718jTylNR1siE/Z1Po2l3jkbiLZ7dzUpQGrvcPiHH4v+g+YRUoV
wshAXUyd3Xlhf80GlXHWGLCmHVVSCSa1ihkjw8ptKi0Haox8rPWYW6zTCKnPem07VKcuDxWEafOx
SuL1RRbFxU37HVG+R/nJiu7tzrtl00mDJ1q1Ucq2/8uB+W2Hhq/d7pMn30/yjrRuHgNBvpXaQ02f
f3ePqbwdqOYJ5ZzK3HgmZRrQGcgDiA+7nUkfWi6ERMG3sFoJUd29tdvBvU8OeydFkHE/A9FIf9Gb
rsjLLwFWdhkkE7wQrsF8s6HLECqxGHFe+kmVm89R8N/Xs4xoRLtkjElurxTQ7Tt1NpJoWEndE/yo
9b9YL0iLPcnE1b/0sL3c7cYoQPiEdUdW+acEoLp3Kg6g4WLAjW6kLQsPab512ga8dPD9b5k5NaYm
1CEn7VIyrAoh7ezcH91bJs151mZdk+44IYyEIjDyRveQ0xByWW84rLJJlv8+q5zt9Zq/duKcri9s
BxLJrXYrp6mvsdxLGbOQkIHtXu9xCJONY65B6kAsuRjCK2fVISdaBSTVjXRn3AqNTClcL5OxoJBF
WrZF7PkIkIMX5iSoPUT1Y7s0DrulJel20GvtdE4VtG43ep1AHTha3Hqo9zbFZb79/70X8ujwcbmK
oUQQqvwBGEiwbMxaXuuDyULGJVatD/Zzoqax6f2D4nL7o0gx1g41JUmRVkVytyMHoL7G3bDWKwQm
u70YJXGDPlz/LixG5pbGFq1/xswKHMAXY3xzVA44cI3YzPDrv4SmGcHTdFnj2m3jxLV3XTgoLN3j
GwJbuB6FYrVmPmjDMU8GtohO4ruKJw7tKCH/CbEKQRqu7zYOzy5Xb4/ZiRkNioibl1NwKj5RKQcV
VBLE308JH80CvUkbeKOs0IElZohwu3MQ2K6ke889ml1IjoV9Q08MqsPzwtuuowWJRDd2ZIMs/mDk
UDOopKgr2Md02NG2avZw0DmUoxjnxzOq6kpxVifl8auP2v7Yd6vm+JYhRq0SEWoJgTW9xjlCY838
xn+c9+GR9OGBJ5DT07rO6nBEApSuidShKNzSKZ0yYLqj2jem81mtfaZW+z0UKr+glA4n3HbkUknA
/mUsomFFUxBxEEVDsk0zQPAuBpQxY/u8gCO1YQnxx9vlC7D5dh93d5RL9ttCsOoOgCVsEWVx8NcH
v0sMVOUG9ZILh7GjmY+6IIppIVvS0S5E2nBmhP7rwTwXIWQSn50iudBvvwyzUz7KDJ9UMb4+b6ea
J+RA+waamOrycbxxKKUZIdFkrzuP77HxJCV51Nx4KnmQOV9H1YLLkbwAA7BR0ROe5G1oBmB6XqFy
oyePVhsquWaX/npiGmohMMg6V7r1RcnblP9/JxE4+HKvGicVQzNy9CI44DIfnTonjmo6V2jjp9UI
0VlKhLW3h5HJ+pbCehsnpjHhY6fsWEDiNYkb1evTMXLuK9ns0kejpmm1v8rcyXAcT2pOguGaxXfX
HVI9UobyuIrrn+fny9lUzzPt0E3p38hrW/lFhALvmBUCM+s3NA1AJWu1yqG3NEXJP7Nd684dch4H
ZRLCJ9Ktv3oLKI38fAph+6tHdExbLFxwAdY5Mze9DIEZqrpQAicAo0bpqZcbBRJpSwITWGinXiOI
KYttZIJD9rvQ84eRTf/wV/QaRTiciNSY6/glMXbgddI2/9Q7JO+8ore02ffxp/7TkAHx7LJcQ7po
sW8b+9P4vOSVNSFBvyrN5SxrlvI61JeAaEuObGqBUhu0X743md2z4NXcmTTY3AHZSq+ksO7Agj4F
+xhXMwie9b0AyLRYP2SYcZ7FzmgXlbFdrHdYujLep4KuZ1Bk8sYujM/xlJ/mijTg8JjFGN3FsgG1
jkUL5FXgF0cUkwwVANifImJ9Ym5EQ/FVQ+HYKpEScHH7wxftRvgXPRrVoJaF8Tm1rGXIHKqt8l0q
muuQJgz+QEXZ//uGHHcXoqgn6hFnmJ6/Mac6O04p4drfzxhsmLj8xg+Z2hQq7BXb9ckyq/N8BQQm
qAAe54ZYj0mLMjZTyIiRWAm/trHhiKuc2s8m6a+6m3lKcyO0rNbYsaaV6qL3ghSo18XWkhySCKfX
XtJLr94854IjSrHTpbrl/8GzKb4xOQVzEx0NomokJvlqe9V9y8XgK7m/rJyzxR5ph1OJPXM5TE0A
wqhqDztBRMs+AKgMhYuvqlMppWIct/Snaxgq9ffSu1TKUMqlWKbVHWiS5Ge1KL5DMwVMa+yRDEuw
91z6JWODpzZQP92vcQif8KEH+Tesjxg8T3vKyb0uy5II8VEwoFuqkL192wab4+rZzb1d8iLyxX0Y
uR0FzlEvNRc9osp2NcbfWLurMvLuaPCShsRZdEK9WpDenfjO0ugcoMCHmkzcWV4lK2r8xIsZigYB
vIR59af/Rk1O3s68heQ4VIlTFeI/iI4wyKEB1u2SrJ7AcpvJ5uU9O3K+7lfAMl5w+96SH+uC4k1V
7Mk4WSsPydetMXjy5B6bI+dRHfPdNNA305pOU0Xk8a1JcM9dYsDvSF8rsmbkHqFaFGOy5qdCYJGI
1GCj3Rs9ZMr0FNUpos+fEWysapfCFgWqQ7mNmUtWzB2VCRsjbzp4oFzmURKzm0FMyGOxT63Whh+m
e7iBC5FYzGoMAi0DFdhUjrEOaNIMliYaDqaEZgjRDPSh86T9GdZHPNpu57y9y08S6xowgFWnmRAy
fnhAYnEYlEm5ed9yLmbvGct6hXDVImu7H8JkXXTj3q6E9+cWCIiieh60+PRHhD9oGSfUhq8zTZmo
DAtIg7zWfYG+BHzHH4HN+zM/t8+S1xwiyzkV9Ijv4va3R9viUV7PWEu30kvRmJJwYESFBPW4jplb
ra0GDVpeycPFeXtvYbVwkzZNuDxmSZl8hlCuHvqEEu4KKOQ4nCMctbp5L8CJJ1cNbtDWMMiq2/cf
Fe9vZynmKXoZtCZlUzzIg6mYq0Sl3xUh4JzxEohKguvpfJkpG1Blz8EUD+4zTbQjPqR0LTrks+eb
MWYGoOjUC0oxvq/ZVgJwI1le3qLJSGwATHN6dIxaSHXeVvihWIdLkDddMeUVElYglCHmJkVSVYeW
YnxGeUNykqJgDZsgtHGCIlf0/nnH0JRpOz7N+2Xas6e/E8XBt0JqLLPJpXwtzLiDT5wQ7eqbMVT1
ln7icKNNPi61AbrtHgnpMjKnqqwJWKMEDc2faqOFzWrzfoP5MOhShe7Cir0C7c9+tPPgoL51CKhZ
2OEkxEG5Na1zpkCbcfg2QJxi1pV8wu0L5NYvMvrlFDSZiZ1Xk3gn+o9+5Q76e8Pwj2KYld+qR2hq
PcAdqggR4Z1urv2aiH9bludAdzOwOWCvrAgs64SZ6jxrxeb6gt+N77Buyi6TdavKhoANIDZD9JGA
7SXDTldAd0gKEvPPL+/4BuS+pMT+TupO7vx+cs8g2O/gDySY3cy8SeAHpx7wqlBsaCDfqvlziKZr
NBc2M3XVehsi9QjUy2nuoCBs9D1Bsu1kVfkhX/uwBHs0pn8mPlh72HAcSNMO52vQfPUyR/BngUhg
zm7T4yyeiyekXmyZOtB/Npo82eEtNhLiQVKQ+Hwf3jkffY3Iq3KgKVwGd5PkWTeY5u+GZK0maCYp
ZMKW1PuW+7ZrDEgV/jbGEFCPQ5zpDM5+tE11RPqPQoiV7JzImUo+x7bfQbqFZqt0kAbT29Q5Ctv2
JA60X4r8va5pGqTqUNRGIyg2Nx01ctizcAEUQCt+VbKrkfTosmF+QyCGANJYJBtr8Ctd+wA0BHZP
xq0mxDxT+x0IcZMB+rvE7mQIE03bYBqQ/Wr3JLEn5oCOlkvATKf4WAmoA8gDhQtPlsyyvvoxzCj3
Hr6FgHuNhY+U/Fi9VreyjAQMNl1wVPESnUFvBX3ORv2Nr8R03U2XR9N3go+SSlAMOp5snzU00mTf
Ul6puYzlRvcSTF3kB1fcPquKJTN9OTwIFWA7NQqvaBIs5kz1lmsE+uviflhfZYQ1W4jPcoX2/nXN
TcngEzFbQcR5kAWlaB1/4NeIDduuwIdAQEJ9sOfqTK//bb7ZiMQElEZcIk0GVTaIL3BrCWKAaxEI
Syqoh9Mi29dZBsSx9I6Fdq+WwX2FcxxkRNgmBRxV71dRub7VaHXqkf2VV3hvHla5X9PDqFgtZ57v
vPsUZHj3PnC1khNCyCE7YiGJ8eA9z0cwJuIiHr72lA0Ic8v6UMluPO3q3AUeBnVTr5OhfrltSGFq
Ypg9wU5eJOZWNaS4DZIfp4jPy5iEo1sypgURotiRk2jYe7kwPNA005lbzfZ+tb9KWHUOFSr3nbza
pnnQaZR7eOxD2IAoIctsL7NM3Jk3nXAij+7v306M6HV+eE0czd+uRYqufDiRs36sK2EiePC3Nk2v
+1tZLfIj7E4eBiLPjSuiTorWpdt+VVRu/P6vvektm8982I/3Wqb1oEjyPkHgVxf8Rkj4VJAd+6oV
bCozl/wq8+6viskYiX3k32FEegOvgh1dpurW0SRj17BJH+CAZXmRJP56uQF48MsJ6REuuwBlFdV+
aDd/097+qBJPiFyKY/xf0WuVf04FfaOWoC6MAOvoMd6VDhXANBoJlz2j1vdwQg6mEhXBrqOc1PRZ
2KDMGH/K7G5OH3FSmsEMF3xsDyHCy3lB7zSA6pNr8ThVsh0WWiV3ueWDYAyb/InthryCxyGIOlsW
TRagWkRxKWD+mM5zPgpAbnrq44KPx4XmjzHTJTaBjaSC3Vjd6Y6s+YB8ksaCjMLZFNJyl1AjZfoC
bwgcqcN/JS1QPJ0edpQmG40IzDt/tyqtxtF5Sxf2tSP1SqInAMj3puQkyba8w8pJ5x5xE2vATBaV
qxqcD9VH/RolW7oZ4Qz7pbfwzX8UKz6ToEQvG17UiTLN3sVttcLHG9KyjVcbKyklK68eLZDAwiXP
z5mwA33uTlnUc4QIhs3L7j14F6a5gMqj3F3GMYkK33JL3UC6CJFZtOuVJCMUC9EBZ1a/jnQqd/lU
gqDrQvDAXI8igKYxL6iwsoSCcFYhHnN43XsWE7ZNcPDhKV7j7hz5USlUimurLEqHZbQGuFLJYZeU
2OSTIqhzf2/jcPCbWxH672gUifye6ds5+2cuNTBoKhI0gPPtYpdbXaMOb+MsCQbobLFRpS1ICZSf
kOcOVSExcvuh7Y1ETol3B9dy2ZbGzaBjJ3ixutrCQzwAa6Ztzc6VWmUmutFzDaD8kYiAlEjC4YoQ
b6PI8z2AwehfttRN9UNKIX4NH6fC2iL2dAUSGAhfXjam1HtLi9DNtTilbgbUnMIjD4rmpT4GRz2j
Cqg4FO6qceq2s+q68y84NI+hE6uacr49bsmyhctQO5sC7bi3zVz55dCel2eF0lQcBuYnhqHzrUp7
LzBtWhBQaa7HBh03rMxE/jqnXSJ6Xn8X+yBY1QVtFGuf+9g6oG1KDRU+pXHgLX5ayAMAsS4HdQId
epV/WI9J6tqu3wx1O2m/aP5gJ1Gl0/XJJIA+1QEdEJyGwN4Zw7q8FnFkR1dhaGAptCwDExG1MrZ0
g6jq4YSMoyxreJmcjMWgGioedQC7K3Fpz1OpgjANMx1VdZi7zkmwNHUJ3rWwriItxkMRUoruYcaq
4SO0LohgPTGhaUBYq9C6LsfZEEffnG0j4b3+kZJS9peGlDyDTVOXNuN1d56/YtQAupnNE0SklGRC
OXr5S8J8vpujAWahEthLVe6iRLJAL2jBjY37cPVlDFbLkmZSXblF3gf+TYC0BBlnt6f8XBiOOBRv
UE/O17uk9mV6lziBFIguvuQlUQtoj2+7jCvCkyQIyJAJ76d+LIYVjF2qrKL/EcoaZM2og2XeJ4Bn
MgUczDYeWsPH0t3bPmcYb5/72l6d4YqCXUgQACL670H9V4vOHxKiRFqOvlYu++C2jOj3BHdm5032
WSoHXoi1ts4ArzWDNGbiWiw3wjHU2fr+SSNoyBt/1emcfq2R+AUj3YCwl5dUCakPmIm+7U6knf2x
jqt5EPpCvajpdhcoymUCV0xkot7oPc0R80Cn2Wc14F5DsjjhWrUahjVcOCurPkuz5HaOM5u+/UqL
1qLxlV4+sHrmDP1K0CwJ620eZ5US70jDmgdSg53BdBs666OkRwkVPWL1otwA1qNYeYZaXWcDPg3V
6vwaFRkpC9m+PY6BA7gb36T3nBgAL8cTCCakW5UT+YOOkSyYQOQfqTpYKNNJNFQ8+9fb/wmu012C
QTqVr78jSo4I2cqn5T0YoptM0caEI+GE/n/yPGmxKiFgqK47Ocls+9W3C0rK1+BrT0SDlDEd1of9
MtkjeBDCYARgB0YpTCJ4d1EC9kVUcbTCHoSBlAjHDEkjJNsv0o1PQKNYZDwr7/LBN0oaAR4Tp32g
rmfI0bILo6TMJAc+NJmqSzbr8PDquDjiNpVdAYjpROLlkuRhoZGBWCameGWmirNF5x15eHwmfbyi
Hgikq4h6vkVQATyg/H2CW8i0r/Y3fBw2vJmohqUh1vk22nR+rzSCmxgBJCK3iGDdT7C+3RaAtJJ4
q1t4t7XpHEFz404tuDaljp/bwx8KYVO1wx/dI8B9WwfQoekrE/Q50MxcjBgWI9pBgp0858Bu6uac
G//6NtOEzqidNwz9xWYO4KKg90807XsQxHuyFp92RrzIQSTBCNGZhlk3BECfcypwzBaK8C3YwE2x
cuu2tBb6Zj7+d3Ea4iJ8YLg48XwP1vh5nCI9rPy34r0YUVIK+EbU9RP4DY02dF9fQMysLmpQfOgK
0iVjeDZ43MmHDl9PMtYeIdjVcKCCpIa9ERlncnvR63QyobLv7FaGzU/EL/N0zTBoEmsmkVZxoyxf
/Fw5PX7x4fIuXGyK8IDPrJDPNVxhVbAVM8WSKP8IVcdEQaDfyXBvQCT8cjqpXowhP4rw8WV+jGQP
m6elI1rneEb6V71FzUJAn75VcMzmDOcMYCI+nnVte56pZaC99rqNMiQen7LdxF6HDqyyu/hLPJa7
ndr9pBRVfWHB8IFzzwGemybQv8C0BDLv9WIM3m6A5IF9zQGkzB68pSri+qdMNaBNki0jnJUBkEGf
L4dmDZ4Zte0az0j6Usboa4ECsIaG0/sRG0Xq/Rtr1wmcUMv4LZUBFh/yF5qmVLjkc/omHinbmUWe
M4U47Msz7QgqrEw69rNhMfke9XmtXIcDlN9ZSbMKgn4DXW1kvpfQxMVwtM3jskW1yFfze2BJiE5g
J6Fs+/Qu1H7ro6DSAf50CJ5VG/+t23GK07z7YVLPBGuiGJCzzHyJaHcvtwvXt8abw6yxQObtR1Lv
o9CWJDZ8UqkQaEKWnB9PkdH/C1+HZ8HX1jaN9MmNH2XxpLPxELC4jfH4FFBV1seI1YmkRr/NUVil
l2OdZeU0rRifcFfauaXxBFObm9vKFVlAFMBd796db+lR5PlHdsEAsM9Nr50dvECfL/kaFWtdvQif
fTCV8J/Kcd4DBkGZQpgpY1uTRDgUlH5s5rgFNKLFeKq4fCQ3SoBlfXl+32H9uBKlJBwxR4ZzAaIw
UKXNd42rFZ+y7/rw9CfhCNKSoGaj3F7SKgm4mOAifvvFIw90oWcPF+tmZigxU0+9asUL4axt0n96
rXRngFkLN19vIqNb/3nYnDBM2I22BK/RW7dKIOfK2Yk7VPXI8Z5hPwrN/NV3fYnWb7qgFcyIYANY
tynDdemDAvRK/w46u4/qhWhE5dWkqpr7Icw5Aoe++8/f+CN0CDuW1KpaKm2Qqf9C2Hyc/oW1s2u1
vf1dwAdEXbPqzB3k4JrU3krZ0shF83hjyXjOQnUoX6AgfKg7MUizkfGq1/VNgpJSVhYzqHybAnPv
ucs90Z/95BauYYCd9pD924W82PmeWAx25OrOSXa1pI7ZeeOLs07icjM67cHueYMyp0/wWqlOKswo
rEr5yeIkwS8RohXHxeeG3K3OYwzwSnrzEtO3tBEmDag4xcavw4u/Ybuhjsb2WnX6zukIP7cLWS0Z
ayntzni/PvH8hOUzwpFGp6RvPUwJXyAe5j6f4XUh/RS+LaLbVhIeOXjf3onSiznIAYqjv0yb5ASx
4PYcBkK6zqKaQeG2jh5dkQJyuKSU9W8Ti7H3+BPVnX6TbWyxW/KpDt2F6z7VvLhPmUicIcnQYfZ+
jtW6AJuDXHov4oQ86gzRogdsMt1rMLW6q6hDgmBsvQ/bGU5QjUOUkeDSB3/UeLukNlBpXvKRo/YF
wQKAiUo7PheiIsEZsNXC1273U6qUR7UlnSr18e1+A8KbEM3dt5jKK/2NBHOYnQ+TJT8sKQAsxKYk
LB5VhTYOFq2NJ2d25C6ALBGP/o8WxIdZHnIgESnvVZN43oUWqX5kqBwb68qXxHKg5DQGaIW1K0jV
gdswATlYEr/C7nMxesarfJh9uayZzOYqhZquDmglZzqVFJvHNfDCcWbjqX4JpCkMJ/mpmHhALRO+
NYOqC3VMtTPGLXTrSXmdZ7w89sSvYCY3K3ojSPcL+/TkUQbdMHvUIpaIMFLuZaolk0v6A4nLntZ1
3/h9bhssG0ycbH+tcbQ3e3djU+XpWKcllE4CZ3tfmzN3QQy0iG570CxJkFdYP0hr3iey3Ub99UXs
cQ/XvucAbO0Yzne+FVkqrsZYDKH3TEN4Mac5SjlbSj94Nkc6c3gxJQ+lTrZCDH5MxrWiAakx6tPJ
hbiobm+OmQi2b4HSRKA/GvsjAQAo7+ugJ8vKXaD5i2A87OxZhl8asOWERPqfDSKbSMbuUMB44iuW
Tmq8EkJnym19CZ3MJl+XSJFiYoR2F6/MUyAb7vFXDP62gOHOgf5Y4grTISpdHBqC6JKs1AFot9y7
tSse+3Y2IU1hz3grxy42uKNzb7BQCUxec5R7HHSkXVt2uc5VYN27i4pVmnyUmN76YRzduGp31Oq0
KLfb+/qK31gjJNo/Bj8eN67zfLP/QIHMJLSqTMpan3DN5Z1KY0XJoJUXPGlERoq0yFH3L/pp4OsE
sNrX8fsfmMyqqVMdCNqvu3g8wukQilIYtaslrI7xif0AFMI5r/3VsrZCfQzNcZQQAeeAAyTaF9W9
fjv3Gng+iMT70TtgO4NTbrBGRdPCqtGdXJXZMYiucNoQPR6VLD0aJTDJaQuo8HdZDA5rU5FqiqxF
Dx6UKswPwZBU+sYMk4vVxGvlrt1bBG4Z2X+XwttQ++M+e9jcNsXtg03tfR8n0lgejejMPFpasXjM
Lko0KxAlS8kPwF3PoxOdSkhCMP70dMkN5HA6vvdfSqIJfMzBChP6fXLoegRFNz7bf/rVveJE8hXU
KE7dHDRPSuYVYX3jElxINrrH8fXYlTw+qcnbVYlMSHMKTX5kKuUbRRvzCuVB+CnSJ5ZlphOhaY8b
onI3ZpluT+p1cUYtNwjutcroZF60TjonUZ4Z+plpxvtdowG45YQ8jbyONoAgKfLh4lLpLBxQuzqZ
a5r9Gjl8SZvdajt932vUnEvWZpql2qavaSWeuCUHapjhQ/Ebr9RW20x9TjZq28m4Lc5uSoo99yjo
ZwxPdx+nVnFT9R5a9+rvt6gbNmvCsrsZgi16ROpTnGZsRe7ZuDfbYN7jdY8sk76DlShwtCYRAjOO
QoAlNe+6m0QlW++mB6R7+WpB4OcaM/cQbuzMgkMw3lH4iEarFucLW7k7XSZdWxh/tEyF8XXJxynx
HCQSIG4j8tSwlR+9KraTY5gjXlkntueE+N/Cvsfa1WsN+SfsLO5dYnY73i1Z3qXqNhf4g4F1OZdJ
kGCipnUFfZkcqUl4UJqAe9i8lJWi83gbprmHS+u+ItIXl95wCcyshR9gieNBz6FnbwVgGZRgUhNQ
1gE0bBEkEC0hN7vTH+i/21MnQ6DAOBMpYLFyiS8tQGNnjbbbZ9z68Pa2/MqagNUHK1ZMv4BCvY+M
aaIot9jxvXmh8DlzI47wYCc40MLefoAAgyDg4ytQL/ehdrJxSpTxxiMlz4iMZjGJ8XuaYA+dAIoi
2lCwUHSaAkB3nmo9RAU67caVdhPEJfzcWg7eoIh3ou1gjsADqFFIK+ndOB7MOjoAMV6m0JQrKt8p
MeabJ+clJ1I+e/aOIQJrzUfkSpHGFWrNHpp7PrT0bwiLHd91F7jaRqsC0Kx0JQpHVK1ERhcSZmWe
F2bKcp4+ZBmQHYTh4hZTQU7hIl2ftYnDU+0hip+GMWw59ANVwkj6R7/yp3SQI7AuTno2iWNbfeEa
UWKTLkFrdZOKPAyc0bgu0hnGadTesyJt1M8OHSGWHnjrIVPef0OhISeWC6r/ex0T9Op5Uh4zRqex
UDbba1AAhNUgXqO8p2hbfqirxb0WUmFnwPtupZ28wlenZppCeCx4N8Gdm/1p9GxBxRUFfU0OA3ek
ERAbyr3Zu8R8bvHpA4muph6qgjqc1q9BiU3G3tjuqxxwmswNJ+hxYMLMpbfI+1oVTAE8gT1jX0UP
kQhqud66YLNQ70Pa+0NO23pDW5W2//PcEUJ/7iOGaYKA8B6BtAJ4Bzylw9AgFfAhRtNqTHky+0Ce
wubS5W7ogUwVosSXlRQ7ZEVNXAqoXFpej0c0RGXmKz4WeXR/gvTIFLQs1vMV9oFn/j/wmlseU/TJ
JjTfQpopa9fgqn1fGaSg02foJOqFGlMOBtDVRYhfrVcNSYoVAC1h6H+M4u1wUJodEqrhbBaYZMA3
mKhuKLIfWk+79QCyvePBFVrx8bDA87NBq2KM4FPyWYpasDuzHCSZ2273TRhAMSM5a4okb5vBVmjH
C4n/1oj0MjhLbyhMpSMYCgsJ780Z9pP8yrXOA2c0mdTaET88/7CXXBJvZf1TqMVJGwojFndoUVjo
ngClzJHl0zEhB/5AmBxf+wkrWDxyn3rNfQdqEAHjgovtgz0binKDTdAVsV6eUVgk2fXjAJBfZjXc
xTQ+U95pr36+TxKVh6klQHqJJtb7F3gdZYBezOFLZuGQIwxtGEhnpYh3zQTWuyByxldOuRylok+z
eCcUM2eYjFgrqad5Y3NgJB8tjOlX1/rwXkJ4mrSaU3ganp7zXJ3t/97cljeHzwpdEPAHtpcL1Bov
mZlDtUhwmMV3WPAk9KPbT5s0IT30IYP/n7HSp4WlwqLRR+wYUry1wccbxQzPlnKqgv1bgjzrY2J1
+F5MAgpW9RROFz5wA70wLyfcu/u10hpmhpvAraXOxzUu70qyJFBt4gWdkceBsjTJ1DB4gP90xkST
JBY6kQ7dEnCl/kW9RslmgmOVR5TA7/Woqtb7EPGQAdaSuPBtFQ1/ie5Dg80WsvMww9Qns1/DGiJP
EMwTRQdZCEWT/uiC+b31Wo8t2hkhIWlA9jXPhv2IeZIZ2dMUqosArtJHD490xDWx9DHWzmp0BIyS
4EljVgHa6LO9jP4eq0NN3FotGEo1N4HZg2hybUiFrXoCZKqrEgR/8qr24EiwXJIyfxi74M/bRGVg
URlIWGgIzbDipfOIumOPeZmhNX1CFVG4+p+RZKl+RtajkeHlglRi0RodCRzPD8dalUOsHzm7n5dL
4CfD9sO2hhjuwAKOSPJqKY+xZZoM0lJkl8r+Z2Zlf5/g+IyV1aCfOGaRj68qtSq2LNX8R6gtjmy2
EhKrVe+OF2qsYg9qlPbWtU90213KEqx4k1wl/2uFU0kNjgux7gdbGlCUEhZoS4C5DACHuzxvWgRq
DvqUFPYGjkPDYWQtzkMnK7T6zL7qwkuxH9d68fPnvTNNduk6khyomxthSd6ztmGJj68hGJk7uWKi
kYR2NiJTh8RTO8fSuAn4QUv2UEeCEfAHkrheXltqfgO2/5S1k1ml4tk32D4s9Qg0V/7p7WG4JiEX
lEJJJTzJe2u0eREDvkFpqiBndte4qPSSVLF5J8fiSJPkHqWqvJEc6QKquH7ToEKh4HaH5nEPyvS3
JQ9sERkVucMcFf9WC2wUcJWyaBjoHRfzfPp36TTNsdgqHnNRSBoTmHu5l6TLUcO4dQ3Bt8azsmeQ
q6OBJ6KXPYBJW0w0S0xa80T8l09PUgLPNdkFZ500bMcQzVxfrK1TKaBWjsydUVOJAhT/SJYwq2Lb
KtpPRZUHcT4cXz4wbL+44zvZBsN1l6MRU0RPoCD74aE3CvMDA3yFMlZMulnxrsBEP3V1TwYCBu5S
M4zxSs+kd6Vwy6P0G2pq6yUNJ5yQCqf0yPeKjA0sYCtgkcOfjXrDi6f2/BoiWjL4i0HPnxyjkLGX
Pf/CQmQHUBrCk76Wzxl/vOZSrLiGRvnZLpwuM4bmtp+dAuqkgIDmv9wCSyz7L5xO7PhRgYxC37qI
JYyJ40mV2NWTiH2fa2N2q5CzioRWNSPBt5Pnl5BjfZmels8NYx2FJYEWQ3/q8WCdpORw9v6COZaY
5rVQgakQf9xvukeLDbOByjXLKkF9HTjhWg/iAajayAuxJMj3ae9uFYSRvWHTsr2IaBl0bCNdXLPM
34XHi3LAMTetz6PD9bCeqfQneuPpD0Aawlioh+yggOkwoNGFxHMnPm3LiHAChDGGhQNrmDNZ1USy
l86f/KUlVDAMRnPz1ExRE2TAfll56cB/mM6DlNPjXZ+xiqvTDRkliq0Q7rQp+xbDfP254+7up5xv
aUvZ1cU8Jvi8K4gQEeLaPaXmXmtNkuxTYf5i/YVuTOtXbVZfjcawKZ5sXI2oYNXt8dB1GktJSQtH
KQFRJrpwgbDVD2yZcO6zeBYZzkwEBTv/0ua7fPAwH48iaPYjUu+SBsO0KQMFA2DCZc0zmPyJV0Gi
szc1O3aIJ240ShJ1Qs2jKHR0PLt2d0NVe596sBrssgYtmSQ5So0/5teuE7mk/7jgjXv4t277RBQ9
WE7ydcUYaRez74kFTYXuwW/HBcKMgjAoie5yRWba6jdorqOTQ9fWAhnGzZfmVCjA3pxlEAXPAMLt
CytaJXcsIOTR/NuAV4i6uIP3zXjEP/ve4ojrTqydo6Dsf27O6metOSwDNoUBhO32EJASVtOo/jA6
4WZBHD7tFeLoLUcV2p3AHyMbytzuc75SF0iqpCqGIKIxq99C8D4jGVoNsWmkNktWqxZHbdwF4q1Z
PyqlRn2aMkf7wo+4TjtNSLq7k/BqDh3dgzTNqkFrBYG1+w0X6aol8k6CsthPNgOp9vw7RPbpAytA
/KHQ9/B2FCCdSPJbiTdcXRDv8ogpoG61wIerJzPeidP6ik6xlvy2Vem2AHeWorQgx70EKiXYwWg4
Wdii7GeRWbU+6zYeaBY6pSU4blFnJFvYAhW6Dhqji17JbZAzLpUTxM9LZIBrU8JsRzlZ0SVxJuq4
FTDlxjlDCX+0c8x+lFImw2gVuWklBWtKKjzEMG9oQA+IZSQpw3ymBnfjXVNIK6BCENm+MXgOeByW
VGsGqKFYbyZheadsHOpYDtn3pVCgsy+qcdi4+7di4Ja/UqJRDe6RpS+zGA8uI61oauT5oS3u+Vg8
bq+KWu8YDH7tN2oegF3H4XaOziqLMfLif9sd3AkD2oWlle8ZXQ9+4HYuVXNHeWLnoXV7FvnxMTz6
NJyqjuMIQKKIyU9a1PBUzI3DagHl24dXb9+8DGdYuUVLXXuIRAiGLMPFcQN8/h8kqC1gHs2eXdk9
+gv/ymImqPoVZQa2FWfqOVazG83vBGMrala9vg+9UM4iGiTwm6J2Mc0hge9dgJedZvnBG+XEIka+
bUYqJGsrBedXlZfW22gj8kjNLLS4ndoX/YNWc3E1mpybTkbpz1W49Mu+rE5c2JrLSvuAIP5N8CCQ
E91mSKbf0be+uxI2B9wK9StM5gUumAGjtAuhGvLuU6WF2YxeplZkWvI0z8Yhg+crv73tokgv0Sr+
rNs2pDwWq5ppbO9TsLMJZ3A4PJGNzUJlkv2l5AkMb+KCgHUidihSB4vF/QaPu4Tbp+/GEsqtrVIu
89cn/V07Z/zXQDxNUOjv5EE4HKTKqLkyGD3W1BRdZO7WW9BgKb8mOLEEqbF08W9GbkoIpFvm+auK
jlx4zItSXTp3TMISlQAvCfb0X9zo4wEt6zcLuan4SQXChpNeG975UftNizKC5xZ5JebKPpuyCBqm
KSlIGa+Q8DGxnRlI89HWy1ZwQ8k8lK8eXkeRizh4ReI5S35n8t3lHFcKnZLHyU4/DkCrdYp5ao56
x+ET0Bo5K5JSKCb1MpO0SbMAsWIVv4LhzNM1zbhQWMop1uuTIPAKo3ADzG7DhPbLmqfi3mVOC8jH
UKdufafGTpTQf9wDZN/TfhaBPqXfTc386R+Wb3OsbOD1e9tmFgxWUk3C+Et0wHx8hrdGhWsZ78Ws
weBVCt540lfnFshs72GXxKDjoENuCey3yjRruju9eh+B3pZ4KhqEau1tg+W6vhDiBYOSQdHeXlPp
0TRjrQl7zszlVgUoRX56vOCrH28ZE5PrpZJQtzqorvWSAwrdRsSV3/EiG9D3p9p16sfb7p3zpttL
UwYLXQldx3AG7thYNAuBm6ZFD04537NYLHH+rNg8q/JpACya+9tGSpSX0uNgqG3qtd5dmuhHKL4V
p6OxTVCYEOw3FyYxI2QawUMo5mz/a1Dcwnn1+4y/iD1r69/sPdPTfPqAcar8yAOcLmRzBC8ecr9X
S9paST1pLb9cJ46r84233q49OmDGgIkXZyj9nP7OAVLXr/izhl17wQEWV5RVZCKhhWJCVNhnjxQN
3i7kXCCnCYzdP/WLidAqrjxJYPgKQFRPOQTYe92gs4rD+TfO8IVkO8FOXCxBEz054yWi/PlGtI3i
mh1a1RbenQ7u13Tx3EDBD/0T6LNNQ9aqmBEjpIk6+2UlnjYuEAr7PaHTVweq//4sQcG8zDeLZ8Vj
XLt6sSuxhjO6XIk1A48CyjBr6Pgeo66bJjU5tva5IlMORf641CpjFn/H4tMAlrmOcXKTsdIgCd2H
uOLafCr5HVUh1NTKQFkjYXHoNqNDBZQuJ/jBvIcsh54xElmqMPZ9hupBrPArBpjwOIHK4GRstXui
jeApxNm8EPiN9fkeWRqd5TiEwhoWZ841BBrQva2PsPDMHcayAgqzIv0+9XmgATK7b1QI4/QMn92b
82rqIDbYJ/nJyFBz6XrsE+xahbxNcUicvEJ9jC9h7QCRmUv0voxkgBn+jeYFoG6UK50rOCLqKO1d
6Il4tkwFfo95QmsEKRNP/DtY5YOmxk2JjoTa8z31Qud7d/bp1wYWUwyrvMIE1DpwjAAgp5J4NuCq
/cM2Zwh7RWgzTFusUw13kCqgXC2qzhA/GQ8hDjTK9he3yTaoh9ITKo5hde6qQMsCvZ444EuV7owZ
cD5EdWm6T4zksYAGyYnYXPD0C6tMpGTJ/WQa+mwdvdyI0mm3NseXrOxsLl3vj23KWx2XGb/ihPWf
SksZBTURRPOnQodJyFvPppk8Cv1BeYJ3GndgYXuQa43nIeoaMJpScbWfo5zYJDHfoUiVsXdsxTuw
khiUEzY8iQQ146UJnmnqopPstcK8oK4miHTiMC8soCpBT1DqAaK97o5807OVhj+XiAZxYhSfdxqO
QYCwxSTtWniZbnV9WjZbOrJvEODBTYHB3rBc9U4ai1rJT3f3ASkuFRyKotXtIhZUzUjmFPOGrz3W
QC1KHKERloUrVCeqzMPhTpH+inxWi6MO2VhYbyTcSglGbwhrS3VXNS2ZEHi7UH15QIdAJHpUhx1t
6B49t5KrisCAO/SJgdvylsYxv1erYh+Q4UEKPGSAvKnRTGEOgvGZgg+Bs3Cq3MwfZFZY8oiTbCv/
aYJZlxR2LivyGQMbEFSIUZxjnnYNCRFtlpqpzDxzA5DU92Ap6zcw+NjoHolyay1Ji8ewgeVKXcjH
ZlnDBB7G99RZiJJngqM3sA/3UCv+3TiFxiXZQ8CWap3n+BUvjbl9rmUk9jXwwcQMzLOM7JOW3NRN
Q9vn9Rql4Ayg113BEBJpSYhdYiAgTzrjwWfhN4amER9AQ63u5TAyTcfCoWLQllGVgv3mKVXEx2Yk
sq8GIL9GkHFScbcsOgSN2icFb5HRMuXTbltUqsDBWU/a2U6FOk2vSiYS/aOYw9M8xhHiPg1hp5wt
p6xh863pH8iI5vrLVEoohVsFeQiNsSwp7cfluxPGqj7oO2p0t5oTM/BLyB3GuJw0hS3r+DC1ubK0
kmVIBDkbmWQuiH1faqp2g8y6+8AW8RFNrlKMdfY+WFsBhuVQxq5VaKOBcH9BBT7+ampUFrof9NmQ
Vqxhc7H/elNRwGfIujtSKcfJcAyup5ejWKTSDvOJPMs/+JTbG7s9uJFReLwj6n98mOvDhXorI/8R
Zqg+Z6U6qQsPyNyp4drNDq4Qfl6GPGCxCU2XxVC1FPUWSttpvyHRz8nR4JGvh4RFFeBP8TdmYGmp
O8mvIcXBQf6+d3UrgT+eEWDS89PGKu1/tPvZWbDWAu++FBpmV7wV7QJQNLuKxMWX8ucf+gvldVrA
lLSpVLBitHJvpvTahyKwKy06ytvRwG3NdNT4/XR+ELI5valL2dnwKTGloYO2VeMC8W8Eg4B5B15r
ZQFs4pw7jsKHKHFrnEmflCjr9wmXG58McNv1bJgGUlqlVBITjzEcmyKJympx8Eu2JsHNxwbCTSDX
vP1RekmZuU4cwgq8V8AdZys4tCqFuKWDKo/6YpHpzvsiKWrxHdH1d4pFqRy6Y+Sn5W3YtyrQNRfe
AwpVMnDxNHyV4sJFlNNLCpZ/WiKlVQMBdnIkVub7ELEukZxuX4XlSEsa2GOq/xCeaX2PVZi5a/Gd
emBntksw67XlIZulTFQl1hScnJorMnBb67A02B5FeNVjklEtywr7X2NxTv4Wl1zd3Ciqxzi78/Lx
pSDJtwK3SjQXlDcLBRIoaEQl8MEopMbhUY/Ct34xUxR9n6ATrGACt6kcAocrz769o8CzTRLWI7xH
CTMt4f12doLK4oHGtAGflQYmUXDuh9N0/po5etmStkApgv8GsKJ5O/TMG+BVciqt6ezuK8v/0NCY
UBnP3djEJmfqQ+4Wh0evmNah2COOPprbyYUQq6AJwlytnpQCFT8hnFPWDWoBUSdHfFwhDhpKSxz5
VCknqVBiEjOmy/W8ueq++iqE0m2xAYlCQf8SJoNoQMxVp+nFczxQ30s5oU5WNEkFxaBl3aWuikWZ
p+6Cs1dNwmXb4VdOTY8hrEquJiyzFdyNaBASf+6jnuk9F3tw3zAybpo8a8d1MKWbF0CrZwgA/1EY
1fHau64upYhvCXmGARKcLdU6uuKhV4/1UaoyCMxRIkwfIpcxUvnyaxznymRpfUYavN5zkROcG8CD
cH8gvTy1leoeLCf/QzSdFLhr/YXQIs/iH/EXvkMdwJ9GcWXvXw55c7Nqd9atq2JKBdxIJM+GdGay
CS8eimf04Yos7eR6yBpKoNl+utXVhfURIO9zfOua+bOluJ04qy6dUQtoAToXwTI2Lil6NQd1p2PP
nLwaKWx9O+ZOYi3gtK0CC2wa89anoc5nM9UMW0uCUNAuUwW+yUgGvVzIOPMO09RdOq8/JbxBKZ9q
118YkdXyW77QGpZt7Z/usT08paMjipUTDGJGY7/0QD2BpwqlMpXXcJRF9WRyMDRmD6mw1VuFrHUn
NRIGupVZZddjG1r+ZHGzLgKyTYpjrR6l5POGu6O4PKjXsOPDZjhQlHlJFyRGTk1b09jt2PtjHc2u
XTuRFTt3V1v32Wan0QM6CasQTQylliYn0KydvAPFpzHjATa6hVhEQxUpqwb534uyz4XkQQxSnsI5
W2mRXnbGYGhYe6wGlnjghcOV0uJyjF4ftbauQ8OCjJovdLxLpTnRiUravdbihj7snG99xb+g0BPx
elgpo2fb9QTtKI9AUVHfb5g5REzQH2lOzxylC/E3DFb8j9E8yPamFCc0h4xqEzcEhg7uYDvZUC16
ZBGTqOjS1nVlxrAivkII7enwsVvZTK2gl9C7FuGTk79zqduy39BpVacvbU1qHEKWnAbvl6S2TtTL
nMoKef0kqYJQKbcACge4paBWYgI9Rz9hkdOHGiGOq3OIB5n8NKW4RnjFUKtsUqM1c70/abVSkINS
0MaLvJs8B2dRvb67HiSnFlQ8iOntUEtgO1PVd70ue/FizPEA7SBBSbZ7Jb5xvJln2Fyg8JjjMHr/
UdjJML5v+HXIYqy755lbyIbz/PU1glsYk5N/1MKyNl+gr/e/3VsmADnV3ln11WbOJQsk+2ppGbzN
Q5ElE0VWHpCvwQZxOSBq756KCo2xiHZ4VUlVGqTOGY/pmceMsUgEvKEdsBhv93Tj45JNAE3Jf+yY
tZLoQym/fx89WlnAVlguLsVJWszu85sRM+ZDdFeQhTAwQ47MXzeDWmpsnTJxhRa1wttCazljdRgK
6Oaqj/krf9CpdjC0YQFKk+1eg3AUANUwxsRQox2vOjraj3FN0lguFHCV/Q57Wxs1tEJSxoLvUcjp
f7AhIlW4KFWZ8uj7+wJ+gVwhZ2AOL8BStJDVGZzVqaYS3dxf7OGOpVw5V2jRrmf9KVou2hnVhzmT
4ChG8pbjERxDCvIjcYFYwOQWe3aC1QvmCim4f755+BYUVpYRU2rg4nanyoivwEp6vhMAjlHDjGfv
70i8yG/dgwa80d6hz7bFmajwhDp0xm+TwYAEGSxkQavyjL/dFxpzNpP0hfwNb41K36kxvtlefeyB
DIl5Whk/uAbnUd/4mXJDkQaH2eOEYk/Cw8ZdtTs7V0v8Kh/qKyilY2g7Wi3uhObJ/HClbWHRic6C
aGf0dnS4UVp+UOnYpsLrS3wDb1XHi2WPddP6O4q7xdb5IkscqqkBSkwAMqMxBsD3aMgIM/DXgfmM
7IxBErlBVz4SwU95hZo+i+pTOjeyZnrA5k8rq9aIRO0ZeuQggTp7LyeEtA1nKi3zUraaxajqdkaG
dCMpciGZoSC0MXLsf0lKHCjeFuppgK29f4QmmkW2wHlCoIj03FPHg9Tnq6dvSFS/7NDfx2Fcg71c
FBk/zQ2iSpP1hLGmg6ntiF4s3eMjdzPzTHWeQkGNu4crPE17pNSmQBLzLzBqnTHGGwK29zSNPVVy
dZi/zodmhhZWAVTLjXE74GW3NPvzZjQXydrARum0HF9gULaVSknC4fCJ37GPhqhspAgm5swFO4Id
74hlbK+nJC62lQ2+kTRPGA+oTwkhaJqbMN+Yh2zyExGIOdnIGTlKD690gXErbtez1gaTlPZgsRMv
ohP3tI5iJKBY8nO4T3T8dF0DHfvzyMiBLMUvk6bxPFF8+yNvdiTL6E5E2Ovj6N9Pzy712/rYXeAx
U2Du0x1WvrTAmUIjNVmcHF9oVXZYNcGR0+7G3aAqwpn/fl3PsVNU4lIf+YlzLHWzzvZY8ARk6xTB
HmkVx6kzH/bVlvi6Q9jjlx9tY813aXYc28awGulTTNEmE8ga2nT3RHAsGFwtIiHDLkpPV4yDxbWj
HBZYJaRg+LkYWYbyr6y0A3xqaaZVZEmFVptkZnT7r0O3mIw+9Qvha43kSs6zSNtDq1GrpMQUkePf
/9CFoAqPguBeNI+g8nk+Jl1PHXYh9mZsX/C+HKgChGHGqmJEqU4o8E823tiGMu0UgHVbItnO69b3
wnm8917R8eZWgDvewa3g3JGhQ06zecAGktL4qBUWGkSMbw0y7Bm8cAzvhRaGORhsVoMPdjozu1z5
9VFq3Uaw90KJgxdc03FhWWcTWfrfRsewQAG2XaeBSKv/2JmyGCMcFXOOuAnR721coYrsWhd8ihoj
dlhRtAnsMoEb6GVglii56Akkce98qo2bvP5VEWiqZrnT3bo6D/1e+rEEuyDudQOq70BWwLOIlPJu
nR/VCes+hOVZPzqsI/eN8CoZmaBh5UH6hU+DcXK+v8p4F5yIqNSDswVYK9qO7lr32N5KxBn3nxxB
BvWOJvmaeA7gQHXW/K4Nq2fGo0SM+L2JLLbG95fdbIhLz2tjLD6MkwoWiAyQ0sawnDgJmXBAcUhJ
Tk7WsRjEwGOGrmjaGFBrGtXMo8ZRf9tssWuWEDDqDLDcWSbOwsFl2kWyVETCM/a3zS9Jmk0i84sy
j2fPLu46paZG70CGfRfgFulXfsYwShvxgyAPMUG+QDscf42f8xZi25/scaorv7uvi9af7X05qgxv
7mDCYlecgGJQp2uPrrKInA3Zh2AQhbMYJ2/Aqm62bbg2CFstlQ5cnbCdAVZdVbSlyrSj94bSqQTw
6fK1yrRE9cHLGEbO2FIaU8FEJNqB0Q1N2Ac0zZfnf5FoqCtQzyoSR3p7RxZmStAeCVVgXruTI9no
xFPkZtti3XpMgpWstY9ef6Yuam0cmYmOhj9N0T7r/JY4EOpmcxvmpxK6DjFFO+ZA4YWPsmkwHkLg
Pjxj75b1hfLy7mNzIZPuMUp/yen2ds9cSoi4+iN+0B6fCcJ5ri8aukWWnqcwesU8IUYf6mQMsJI5
jsd+pug+k/jOcquhPJoqoXY33mbQPc+Q5tkw0k1C4poOcAxZ6Lbz0WRhf7raL/DJFs/hRnUhEiCA
KB30c5UXwfSVzgZ/gjWHJ6ZDWCsKz/0IzibjMfL/jGPPbV3KTagQc66i+VKqJ3jzPiPU72doZpTq
jMP3QlanTuomLCgxM02D/+10/34qZ/qGPU8w9JdwTyks3qSmba0Xrzs6T2Jyk+nzy5QtpAfQc2+0
WsAhZA73wS5oXwIuequ9OffLUsejJt3Z1JalTmkIbqe/KdkfAyd65LyWTF7X9Ag+RTOREwWslhbS
GD93u2LNAzvIn2mAfVm2DUaT8Mx56JGxTieXQefiDKA71sRsee3bayAQRgPnZUAmfOFYbxhJsZFq
A2D6s+N+SPriPvy85NgReQFziVIPAO9ZbDgimi29RFHjW6JeGkpN8eBirfRATzRyBFhBJ36x8apn
YsAYb5+XFFRgMaiWkI4MPTZk0ZXtElArmycs94a+vN17pX64qRW2zvnMMQZ2QuM55Qd3Rup1cm41
FTVI4AIQtYpCCaLWSTCQ36Gy9yqNsDWMsKTVubMsV2FrhBp3TJrHz70nCQwHtZvBdXbdgn4xZVIb
EnjiyXcCO8wuezQtVScSHGE+6moV9DjcH42Ep1KAZKbiHnKvPwyT979q/OROPh2SGZ2wNDBEkgAG
y4RGafCteDE9E2yhOAHReWl+u0QiZM/xgZNK/OKW2BCiM5bu6RDxRyAmLQcq7zeqUV70soYFrVjT
pzyuwr65kEtqDU2/28gHpOan8LOmLJRn2y7acimQgEXFowtzAr0JiYVQSxRIOTIwicY59rV17LJE
yA3j5vh0ByMq1UytAh0VIRoX+qJNejNKigczldYIoV/DHdegXW5JRrEn9xOTvZIDHI8bZzR6s5QI
o0/aVwbQMhUr7f84Ep6djJX1yRat1rt3uw6fslkBGeVNHxwIgHNHVZpOTsuBO2rlkmHQ7WXc9z+i
HZrjx1MdQg7YGEKh+OWeBPaIonW65doLsXl6ebaZ7EcicSp1ZgmfnXUpsGKjOeynpgsq3bG/gdEI
DkCHRXfBfm+7pgKUsBRf2NT8MH0ZnFVSepHnnjgIb/1Eb9y0HquFu4VJI1FdYDqJXr6KGec8jG9H
9FBOl3+zXK8tqTCiJChecPMVym1Nb40Qdty2cjrdGc9lXJvoZcaGUqg+HzDg0zXeHUZwFKiy1xoi
SbxY2PTkb2SRlPPfJ+qytv6IQle2vOzM11KgpqJCj/nhr0GM4UvdWtTk+D/FyGJSO2mQkMUl5ZyC
dH8YrFuEepJjyDiyKesFUDYvl9mW6Qw/XaihV67ZJaD2J3rrO3IENmS+sL9p25jBCQEugmrR1Qit
Fuygmy5MTNkdJlvIXnkvB5Zsl2YCdmj8BuSpzvhmyZtldtNW8wEfK6Wu6Fh5SP6jQMMO+KpROpLZ
SMd2VpG1rjc718s7qqcjUK9LKzwb1Zr8iG84b2ZccLMf72Y0ZvNpogHvarE7v/yaegxP0e8kYJCh
ItDIQIepPWAACwMV1T/PR4EMTw3wSrWckU8zycTZ0cfCTu4ZT8mgrWjGavS0IrK+GOeqyaC1Pkal
ChvSF8w9wCN+kHIh5uRWNZLa07+WSZobZwk9cNT+V2c+sq6YgH7+pDao8J7oQ/h2CxLPXs3bCz5C
RPB//h7pu7w07gSZBgzEUOWgK2ywCf5bwR4+O3b/1WWpRkQhnZAFUvOw3B8JqwW8468DxstDiywd
0Gjen6liSxgKkpSZ8OuTYoDbI2QCbs7Jy2xM2QUT7v/dlYufoz34X1cBxLgFTAH7vDEyJp4W235a
V+wVjkG9Lj8XyxyjuCVmF2uXqrQPMSksasT99s9Fz0jYcx5X8UPaachIbhJiJQ80Ah1uTCOoMhZT
r9Qpe8sR6zLbPOSj3fA7XWwNSxq3Bfm7QVVFZ2E2WDKqCxxvJq/7pqttVaOPxbHc3TC51G2kQAaO
AfKGAX5wmopUIzsZ3yySr7y3j6nrqTX17xVTUWl+1jtLEppZrjeuzKJW08DEi3kkSx5OSXgcQe4V
HG8ubY+G0lh5lo0L4QvtZxoWbLAsotur8ndPEmMSCPb7G1+VSmE1nPI0NZqAMlvR3A+Ut2vSgg/U
ZbDPH+f5jVydQhDtrYu/UgmqFdB9jzMXqwGQ3mEBnLmlg9QMC1uT5CHpagGZRULxdqEJWGCx0Gw0
yWIzcUvK62sE9H2QthB8EYbptzg4039g7Q2kYfX8LusWNa3zPRyhZ0SjJRScaL4zG9o1Iq9ADC/J
ZbcynGb4651oyBZ7QSBKJ5Zf45xZeCyfrIUbe0XhXVml1JXvy/pX4d3MTfvk8ShtsxunoncSLDwl
HMhOAsVzjjAlZoBhHeP8P3TUCa2q/u5/oFzkLFrQoOyol61diPZNFq6QCLsraCWbVuSln6QScZl/
gP4Xf9ftkwdjJRPtTEy6D9POgKoxTjXKlGrUGLqdJ7YWGCnJXSAewYv18TG6WuWrY7dSvujOlfMS
XJ9MjGzSR+aDGGbuLBx8JSpfNzwdY+NfxGwi0YSUQBrMbWIAHTWxqR/aWuUm1loDtE8mDETPBpzp
/w9YAZep2CWan99+sBYod5H4eLDa6ydflvZR86KSr/FepH4DD/rXUVpyQ4l4eJfnb8Al2vzyFYZ0
pTTb9neHCfkgt4bXZ0FIu35uTeNpMzoriv6U0x8U1LMDnz/MDmtZX9W1YQvQuly3IwJRkaSVpR7L
wVxd9LH0GTQZpc8EcLwLeW78IEYLIOGRccoaQqEhu33HJFuUhsQ2JBJza2yn0ugH2IKcw95pMHgY
dvJtHK2bV5SKRh95AWBJQk6izUNdcDmXxjH13NOAUBEldcMhIzfFUluCpLrKshnUCdcAVUHC7jB5
XlOwfa/9+NmQ/5XpUBug2xZA8l0vYkaXSfztvLt/RdITwYO3r+JCKnPDY45eylHPxA07VL1REjl5
KdhnvTv1Cx9HsYoDc9pYE+mimpcySK2M9HGb/H01+8C0jmcZgKrhaRDM73xnbwd1VNEuXY1w4h62
1+1ReQQd2hr8my7HxG/cUsyT9y3xVzgxbnx2eezB3zuJSbAJqXDWzsjOLFZwOB5O5t7tnB1+YAjt
S1aMKZoNccSIvlTEsEe7w4ziChDwRP1MmXSSyIf59jbq0GjeZ7LleysgpPhR4LjKwb9hU35YjXQV
wkOD6xF7vTdh0d4krJZQXmwDv/BjyVLc/v8zCTMdhfT0Ysb/5vXlhsAFDbTlN2zn9Vrs7ZpKIBcb
RLwhKSWiU5YRp2bzNE7DO1sVGjillj16maSLWRnMMgC/rq57ni7Ef9Cm2noQRwoeApKU20uRzZ1x
zJ5a7VbhXwWNi3t53Q7TY1aijkF6J8J0dtn70cBUVFqdaqMxevrTDRCFQ7SKFAGKgBDIoY2TVT52
n5RB27KMyndA6te0XgZD457XPV5cAPwkeGhNx1u6MeNoQ2kuh9w0pQMjaPJ3nSTQGwvMzfevun03
3YhsxRMnKfs+cdnQ9NAo+4cz4uqYUZTutGJIR/dlHC9+Bc+JQMyDUW5EO6UbwprA0wq5wpLZL1Pz
qQBUFM4JeswlUzbwg3MKnu3oD0D1WngRjFe6dobBkGAKOdp2ZEHGFCvCCOERLPDE2Gp8U3QRwzM9
w+x3A0SKZ1qEF1eIw7fSobap9HO5RK/TqvmnHJtzJycZNuDuEfHvom4XLf6xcCS/Y7SoVLnjBWzg
2uOMKH8AGpYbBXxdYEBdplgl5GmZv7skjGf/VFu8aKBvIiB56ZpfG4PVOWrmvnN17Fx7BDXThuDZ
hqLJ8E/YNjIgqKFlPQFqvZNeSwqi8BK91dRgEF5c7XeKWgzaEaqyQ7zU4m2YhTtFuTaadMuh3NrL
od5nRk9oKvVTReVHAPlYwWMrVKmaLXkbTdgwbl41cn4ZNQL26GzxIT3r+NUMPY/5BU60qAw2EJAs
QayQYwcJWEJeOG4qUfNQB1vYgEJKsQ0myhjU3Kl09d2lYmQmW0eFcWXDkUFMc48OY/GLsRk+h1z8
2aVdfVp/hy9hGtqaWakgoy/VqKvbsS53b3JjGbdIWWjGo88IQpmJhLDu06ziC/4dZrYjUQDEK3a2
Edm1z0g/lT9id9t2rOUt3YrNeMaZYU7mverFkyJtQUM8Mwq9zk2yKasyCluGUBgukz15dPhsAHai
p4XXxX7ae/EfJgpE9LXyKnTPmQKg50yB7P4U8KlqytNcMEm2R5cWy96d36D7/JuASnLAvKU/FXEf
n/JlZb111msgzFr3ly4T58K03HKvDqgwjl2nCkhdwL4TObr8kyFOh65AVCxSY5vv0EyBqQL3AnSn
72Nd1mM9Ldd/tzlQHYPF2KOeGgFZtra9KByJH7lISnM//WD6VFVRjZsK2NUG6QseghleNpXcxHhZ
6IFjybFQ2ng37906+ARgGvcd3L8U+rBK/ouyRVzvx085A5irgvmcyHKqifqA07M037Gb+6rp7omH
WvNpw+w3YwTMc3LV2UgV7XCcFwzz7DaRaov5XyhaEii0ytzUilYobdb/jpnmZPbhLh5CyoDJjHss
q4Puz9RPiGdR5lPuj/ZcaGzVHLqiwX7aWNkqmUsjYsMCkTahTOrodUTZc4HOL/2mX90Fa4vq0e+3
coYpaEDXofVgIGnejNNIclZx+4tEX6XBszE3WZ9FeiJ1cg0VMPXn7C+Z3faNkcnYc+LL6yHw3KsG
xPpW4sPNGcF4iKXgpxJel2Te50Uo1X+NDl3bV1FAvFjbhl8SZLfjNcMWq414ZOdI0x45RmrD/FT4
uy+nUJMiN7PXjoK/kUmwL2nmiiUNOad2ZA+cz5xXFfCyoUDprvLjUX12i/G5hV/2vo4gQjhZjOH1
ZppQQTFuZlcyLl2vi/VAXlU1zerzvX7ZOHNPKKYnoAfMbof1khJ7Ox3BzjJUwLIbN1N5RBj45hw7
wiirLKgH308LLDKHBF4j+JLFQmYHlhcU4faKkZoSCMDaeJydNkOD7LbuwNkvqnpO+17NsHlBXx+1
mBG3d74toNL1RiawuqwCcBWqmbMYm5+qkjfx2GoSdI8KID6vjsaKDJvVHEyOxj1YynuHe57jRn94
Bmfael2cbJJkySDi3kt36yzWGuyoHW2evoqxc+o9cDLjIvExzF6fb015IGVuFSRE8MAfPhRmHv3n
juIIcy8Ochxuzq/zenLCQ+wNsARGCC913FUrKp3RgAh1YOPr6ENXXzsbk9VSSyk+FtVeD6L9rjTW
55Snu02RcOIZ47BTcRv7V93pd5S/boryeVdPo3iBXjwqbsJGjzzZvMUWDaKqsuUFitWXMdKGhHOg
QrM3cRvfGn0lsV1fmBxJMZ359x/Yc6Sg1zSFfuXwosS1UN7MJQlZr6EXEcdZvot3lc20f4dQh4QC
mOOfmC+q3RsFbhbx7ptcXzkphTkDGbzg19nF2LONCoh4IhNaMoqsQNBFpAkdcdTYO/VIuEqvG0fk
Wwrg/ezajGY0rqTAAOl2Lgig/r1HlMfI4C13ldYfRcOVbg5Kk/8mgdoQ92bfjTkKf1UZ038UK6nt
IydjH40CfG66AXXmq+YP4Uj+fbOhZxg81v22F1pomujZ5u7BCQfzf4Dn52jp5xcJoYWZwYvQoMIx
VESfXkD7nRpHcuX5j7YpuGbZMXsOEiTGh1lH5561YvmVa1s7/zcTEuxLAQnraR9WYV6XCk3jHxSE
FuHObtSe1M8EZqjtjSwYfenfoEXMOnUq4328Wdc+IFyt86IrhzJtN5c3JdhXCPi7O9IBJGKBNGdU
N89iCeWa/n9tA+biElJMntkYGkkOXHP5YSTvoi4awV6ayC3yFecBHxPMwaMles7C5Bro04rKG4QN
k7VWBIXGZv+JfIkfMP7dWgfKADyfrZHsoMVh1+OjT1dxTwaPKuuvvy57JliafpPJuvyT8KPXpSBm
1ComTHi4+y7JuA/H0UkwMuSzJLXDAEYsQ0g5VRvVbJGUrjNUvqRi4nLaVbETiJ93ekBnzDE1qeTI
5hfuAF0loqLZlV5gOxBrLecglaIyOEc2Ywt21T9W1TicGoF0A9yjlxVKjyRxCaipNi+7+UgtNL4Z
0kxM8hzEpBexsIzP0t6t0FNkgS8i6sjwvSLW4oVwdyVbNw7NVrhxgrzv4UGY3aBZbT/EhlTDvbHh
dGVDi9IROkpbm8aihL0kyq1ZImpV1LxuJxRHtWVrGPobOVb4/GJHFmGwrTsIlmzFEDUU9WrKHJh/
TZGJAJopcMf2pQHrkuluqvFYTJT2eYFltfD51cXOWOEUt6+0L4bDsKZRaH5vJs4gGWYkrXbkEnS3
v/jqSRwVcqBesokRCzPPKQAbtPi0G3cV3oJSDc7Nf4nCUJCmDB0Lqr5De6k3PHdE6wTKz0nAAJUG
r3eJO4IO8Yd3ZweJpO16J9t4CE/iZdraAnZpGxzS82QpcijAJ8Pf9U45gpr+Fl0Yrr0QO2xMxvYp
iuU1mJYU6T9apNh6gGnvDMUvbFO41kqDxDY5Ze2vHY3AgCon/PKHFc0LrN7m+34vEUb6wNxOSOE1
hevJRWS3En1HV7gzlzapcEjt1ioDXFRHg8vgsEavi9gZwWPshg0CgSKu/Zn71SA5BfE+RGKWaMSK
hadCA9n3VYSE/fXCRZBnxbBkARCPi05j+XR33XVZMY3VKv/5RKpoEr0tBSc0KJnDGqpSvJzJ5A1A
IaSQLA7VQK6nJwmqFSsUnjCtQq/oEuOsZHbptO1D5N7JYZc/WzbXKyNRH870kVo7vRGndjI+yoRn
9b/lB3oNP5id0YvHfWm+LH813Tdyc98PK677ksT3GxkgRIxChEs6cP2pycAEURsiZi3ENmFBwZCT
FlxTMbC2HZ07xe7894Yq9h2orTAe0PdxO/9BukxiNediE/pA31qwZoF0aIrAnmgTuOsECOaPZ3k5
uaybKpe7ZC91WbeaI+4wqrpw3h7GKWIOQ3b0e2YA/wooipNkzWUqcukm+OmVpLKXCIinACqIoCF1
Mwhb5j01iStb1caWNLEQHZNmvIzC5rloonAUUXXIvmeF3ySLtMG8hC0oUWNnVGC9llBSMAFignnI
aO+DCbtk/ajM7NtVeSKRohocwWGg8Ijq7Y1ldhkVq8IK5AY7iA1sql2zL82I9vtE/iRWAeZ8Z4uu
NDt7F0/ekJEvzMrYBSrjYTAVe0iW4Py9u/Wm/L/kErObnWY2feCtJLDF6IknpfCDUSvnEl7tX5j8
RknRHZgca1nlEr+LRa1jm0NcSY9As/KpejXzovh6VVBTVCePBygkAXmhCuD34/gbTv3UFfEtpxDu
jzy5wALVmaj2VL02QDKXfdyvXSyAIAlKQM72BRCr9twfHeqzl8Xtb3zdSVCkCuAAk8wcxGM4dW4Q
6DGpKzrEJH4b2g1z4pKHzXFVwmuTgkd1myO9cCgJoFHaA8coa1Rd73/IWt/OmB5Nb0gJ809lLyju
WGlOuQvHCIj3nU2g/9SyCDJyWhc9p2v1zoPMeWWIX9ny3knmz4Fov+or1KU4pIWW8S0Kj5ZihIRR
zj27LE97fUlHz84bJ3JsDeFrfjLu4m8KV9P8QM+ZqFT6RE7ag2wsV5gWFZJwdH9bzpXqd6bgXr08
dsyuE5gehrZ2V0MWz0nL9kee/DZxwlHvsiAjRlNuUKgtIACjcNJ5GBqAU3f9/R1p7qI7R1f5s4vc
Mky8SRnPe26epWHqIUR8s/3ToQQqUf4ORc0nWefbKXioXYiTCzW//f6CkWkGTLEauOzAHzvLFOvr
qrjaUSuuY8nAwW3WLKMK7PvSYV1tzavnrUAeZOCtOi7WV2pEiEq8PeCDQUFPPFjK5VqWTJQuH6K7
t4alKKs0b4Yho5zcFQmSFs2578UH0tiZn1S+6ZY9cNLRe+4pmCLJW3pSMNL49/dF0qaPRKEQWKKf
KKUtyRJgzKOD/ru6eYTmsW92sr1HNtvA37v7ARSin6AXjJDsFcJKa1bhE5tsiBHdCPdvUbfjbx8V
u/Xha5Qc4nExPxopCxeHPuLaHNqGMNJCAf84kR/MnRnBiFmIQIis7S0hetaBtiOZFgXZoFJCqtLz
MuEnlheI4XPnEYhmZFMSxw44p3aK7EX5K613FH+K3VtYqQz8b3VQIe56InN3CuHdqiWvrA0A7BVY
zi4nEdqeRpu5Jy6zX6sUBp49gA5AaWnzt52acWd4DN2UHQhwW4O66aiwStsIi+i7ZwL08rWx2xZm
rJRXvG2pff+UtpB3BEZIBLXf6ncijvSfU/323yAVV3JODECfgq9LG461DkClCfAVGE5WZY9I6t7B
FAA9LYiWCpKsKRl1v12EK6wazM5G6cuD+s79NNidSG5D7vQFkjVlx+czZbOCFiDhbgVZnFzy2kD7
Jn1Pj8X2/tvkOh92QFPqcJdDPU/PJPe/Epg7DkT5mZHmhRFkTePLCD9a+w74HQ5nXA4ugKXcx+17
JrplDJ+IHLsHyJMhsl1BZA9bk6tYzqZ6XIF8vTNggKwqjWow+h1pE2D6717ip2iPHlCQm81gMTd0
7gfPu2yhS9XM80IdsBJg0rB6CsLcq0UD2UWYbbYKdA60Lbq2wlCAu6QHwTQlik2WunX6JZ1dOTpB
6fu8MrCEfH/hiwmL8QVdjReYpI4ZmmbJTlV1YDaqO3njSZqBexGBVuY0NMTqw29eOCAOSTBPxxgS
iaPnLn3ZlRpeAZkOAKvupeTn3vLbSr1zcL4lF78EP/109kh/fglOPzXudgPnxpyHPnQmJGviNvZE
9tHGNZYXNoxqeZ/5NMVfKrNNrHERJQbAQJ6iAbtoux4A7qxQqbCKfb/lOWnZklFmJVsilhIR+01A
j1KnI+5w8eHxHEeQuHpULU3n8laBUlFmtGruCmdcGLUfHdAxE0eHVmmNXR1Tdh6kqXxVR5jd1oyI
SrdfBbEcpK3yru7N0NbWWr5bAsOcN/8BLqholVBOqDo3/U5qO4xYLTcSsG3fBtFKJzz60V+mN4/v
6SLUWCQ0kimUy5PXN4U6zEFPxnNp0sVyqhRQbIjJaB/HHBvRVVbpOeDBwmovP9absgaBhw93GDU7
XBz2Jly4W0rhzvSDaAZAylbRz38Wg58sPb1Ogn+muBVfRIrWleCPo0iauMfPe+TEa0TlhhihzmOj
AdRUutyiJfo3BJrSOAinJQF0OQj+72xmoOv8WvKZ30DW6uVlOq7fF55kSUKTsU2W9pgEQcMhidcJ
6zblb8QGh3bTwNB5Q15sHSDBVbvaOLBRpPwe3J28ZCe9Vpn28Se6Cjwag3xkEcu3hVerJOw2UocI
xLW5g1cFU4CsXo/1/k8G7BbcbTviG8deYFAZ58zfJkNPvr03gBazg7ikIrB1zP5gPbNjSA8lH0DF
xFrI3mHZmJj+Tz5AYOyAC/4wsPYgUlWFQ6OPZCry0moyjFv5fXNwbF8i7aH+MdgcUHCLkWzYgosa
gQRIuzhFGd1WovczfJeI0o9KC8TYwWh15bjzLBSHfY0ASuAtiQvr5srnK5F/vryc4gdHlEKwv506
21VN1u6m3DrS0pDk0SDQV8ruaWTBN/M7ys/ZcNkyjkBWnulIxLELj2EIlO8D9kFeCuKNYuDffupY
JnLCo4fmATvWP8TM36SGSsln0xdIJvwqGVkTlV+7Y8q1xI1akKjosGA4W/te1y7bpVmqs8OMk964
GSWaEChfN4AKLFNMvS1UdOwnnUUO+E/BG45DvVjCY21JMG7FIkN4rzcf/KY33lt+nERFds8kCdxi
AO8ypw7fofhxbLx3Q5Wcv05KydGKRTHKtuvj+adjCphZOxQHqAkHuzFpWIw2sZ3v+bKbr1qQaNlF
M3td/qtXhWN67pgmDnaZqN5skRUun20KVRD9wFF8bCr5f8nP0UzV9S83AN/wRRy5tDavzgHaItN7
kSUbk5h5gkXuAYCoXC1js1gKkr30HgbXj+KEf9qWsQ9j8e896BKTc4GXT4R1oyMn2wBxrxv4tCV9
fhiboaqaBPp1XkL3LgEhJwdNCdaY9g50rGO65eNHgJesv9euOhO3NGRq/I8+bPYvOTlb4Q4msvNR
0fA/b/1u4QhjNK6+5gfTYxVRYAI/96a98awkf7ECDqX20J8zU1xJecoPDhCxCHYgaISE97StU3QC
0O0w5vvOj4ZVx8IcmHxZ7uvgKxzxtgp1VgombiAFCBjql+sywGEMsARW2nvFRRXozmJAuO/g0U4U
+doYJbzVaS1LE+8wPGyyEgGqVEF4M7vlV+frzDM2CU5vl16qSOc4m58+gPqv8W+PCQEz0V0dupS8
eGlLUCHYyeZLSyqbHzAU8NeWY1+ymHYWsGTgJ7k4vuon5BVI6UqWanUxQ6q3uWLE9avZ2GpQDTAz
eM3x5stEc+QYw3FATwn4HldKKUdYY1bRIegWx8GbctQe8Ud8RXntHWzMymN2QYk7me5rV4xSRDIK
HSoDidIAJtoxgiykCS1FWdrqEskjNZtCDY3MOaLqkDhkkpBp9qMbQSXu2FX9b6LtrEeTMyaXGN7v
KM9yAqRLzsw+9gVqBdqjRYImjgiXoXvzn5XJLeCJvnf+e/fdPCNZ88Um5F/FVj5eThITNLek4YBs
N5JrVqFTizNOgg1EFXQXkmrNz7Yj20u/GJzPvaYb0AQkuFavw325ZuCzPREtl09hGIH1dvWf6ODz
GZlGroTISnA8uyGMiKQCOeGsniDBSj540nyO20oOLb/4YTd28YBUZjoxgR83Ug5Vi4tc8kyi2Yeg
b+inPrdymau86fVlZMebgND4pOiqhsIse8W7lS8q8EVrs8Z5/gd4i+rt6QY9fcUAFrYHTBFapSwO
Rh6Bd9W5mQL9qyW/VjsEkUPyvFwQ96hHQA/4BcNtusomBSn+7zX0pkP7iSSd/jlx6fxMsciy4/ew
Y3JdAcJTSZNKnFUNp7DwaFWqU5qUKvSsVDF2MBbas0jZaFvVUBs45TI6MryujvpSi4js4AQV3ewV
SewlIuiBL8RUYuGvhKQqxUv3M13Ysato7wFqP4aF7E53EwxKYzh03/vc10dNBMiSpFVb0CkdEg9O
gqXmFQVbcAHKFGXQrrnRxBFs7N+yvizYHY+ISvtsJTmxJUsR8eJyUTxcapSUTcriq2wuwkjhGJqs
pt2f9TyN3IUPUqGyCkM9ISBspbIXcjXaBdpsFskM/UtRc4bfeNtysqBE6MMujedqcA9HiFtjkwdK
tMgXPtBAdkdTwC+6BTQ1XULkQZaTtg6hKO7oMZ6G0wrxfrs/LVta5MEEWKlQrp8/Ulp9LJoYijUt
IIKX5z11950XalgqkdsGr/YOPZYsaO7UiNC9/s8tKcVP3torfEtefTBNCnSeTQkCjYHWeKRcY5FR
yuS7wPT7ZQI0aXBCAuHjKU8BY4X2SGTKZhDb9fONUp9rgmySSWMHrVZ59OcMCpanpLTll5VsNesq
iXDuVuLV/7O72/2Rys9AUMGScSliztOgf56IhyW34eiwkP8c5vQzdToh6ZpiFrIeSfH5/SE/+s2w
5dZfjANW2Tb3QRAVnFwci5rs4QbUIa5duwDn/TMOWsykjuvCkBNNZozPVFApkrZKJWaWjD51B8hK
1bY2z8gtmM8KUN4q5qEQquMA7OZOme4mDDO74c+tNoojzxyFO8MVkAZxCbFEehf3ElAJ65y8ANsu
s9gqR4Xp7Bzv1fG3GUAsTEKWNLyZRG562ocPpwXgQ02d+t8MMiJ/RhoGv9pTxECJWW6SNSwhYFeG
HoPd6wQEfT+DwQkdr4osyZcUoCUDGxO5oE8joVlJixeHdIhVXFoEN044PWVkHtsNPWr3atvWB0DY
awHa6AeTYPWxRZMQCXJoF/SuR0LQ7JTmI2DRCQBGjtrMp2vhB1AjnWTKQsbqrV59FMNAO5tuvZ1p
GW+dYx9PXT26KP8wzjKgXO/gakjXpvrgGPf2Kedf1nxi8NCJsLmJjuh8o7RNFP2/8qwxI20PRh6r
u8PgA8dy0ZXGab62d7feEjKlsw/1Z3kfcwkmhjByVHg7HEWIxJ+zx8j/ku0WvFjBoZTuwyDhehBZ
jKV38LJUdU4t9GZOG6mmV2IIBQYzx8YB50Qs9fxKAngoQM1IqO9BVng8fhVgXCLG72PtRHTNAlBJ
/24+obGA1wKL5iObv7sFl/D8pOP3XTicpNI22ONd/LbS+2z2+nlDlougrdtFTVFW4+Cfkl9LIhZj
IdZojlF+4da5W8djxxS7aDylqDmCe7KI/OB4now4Oqlxc5HXQiy7tNA0iwwdTs9UNq2YLm/j63n7
TmRQVyNOfk93vQZJpl0tri7jW7z4w1Lms5DjJZ4rhLZvhXuL6BFXi7H2RkezReBB/Ri24hjCVDqq
T9wchNyWi5fMi52r4y2KLcrc0iu4owt9m5eesuA6dNAoUqG4eSBXX9NAN6UsYt4ATZxJibDFrBvr
JBVJtB2AN8w4pXfP90ccfmY/97IrgHa6tiK0Ebz2xJNnucjWFcUFvCfoMT48WpO55GyiJTlImOej
a2UuqxUgl3N+e2rmNXBCeH0cRp6eEVP9QkeUkndrJk/3Bm33TgOoGk1y/1r1E9Lh0tfG3eOQO9uW
naq5Mej6QtT9lXSmp+E4tmNFdHCu+LB7HVUBTxuzrwSR0YMkbGtNQ7hmZwdhS7BOjPV/wt9lcIeC
2OW671DBYcOavL9Hi6eFSbQTExVfwutn1CUACDVkt9/XQuVBqBRYOZ+Mqt7BCxEMnF4KlvDrmmg9
MioYnJ/lCnGnh+jNYfgNHBYBgjPumPPKD5ZZQYLttoQEJMkcICT0ReuwIPToBqPdCQhLlrzH1UF1
ubYGhFgH/pk1f7JL/LzHDdjZR9J1B/M2QmRqbyLN22ka0XApTvnpcnRQykl19whKXVqdaMZiMxXo
SiVo6VTKYzPJu/QxBgusfJ/1iCMm2bTMRu23vwk/AZEw0CXpqf8GULWxYlb+vybxN92bJm2yLJ5j
4jb5tOQ/Qhd73lVhJaDAna6MpItSdWOgs9n0fdG5ebHsmKJkdeeeNbXX8u8CueRwiz+jdArfWVk7
oe6+mVGm8144R9Lm8wVl2xeowqYLesL/8J0LiRfoa5OAKUVxcCct6KnNREaAaXLRPaRhmyx4dYP5
BQFd1kyGRktpWyr66duETVtJmOgAWfB1MIvKc0IEJwpye4kadmHT1ta6xE7eLdHmHpSHHN9ZvutU
Al9+D2v+V4I1DE/R7TalV6jZRDYgkqcH/lzc5jcCVUaHldX2EzM/OdcxseYl4BigxqUOgmb87bNu
lfbYzoaFcm8f/ldRsE5MKEx8a5+2DO6Hx4ufFY0okQW6KULziax4rztG5HOe/tys8gpNRNTbsU7b
saBQiZpjWyYtUtJb0cllluggGc/iumlOwrRqJQdLn20K3Fg+JMDtjQeQkPdqtmhBF/BC0lcak0s7
HT+NOV1r0xNoBx/u6pNCr3oicG/KRHxjWLawU7UENAzy8GHRezUfc7JvVK/zc7qNQMM8tMwNDNLG
jClOB7oW8NmFerlgOhx9iNkLQxL5JG5RWzIVfbHAsPOAdcGMXK2WEA/CZPAFJeuE6m99k3Kgt823
YyvqLpI5v1GQfOVOj6vZJi8jiS/dp7obwrcDdJHBWbAPDd4iZ4qj3cLfUNTFSRViiQUfbnZo17ky
QE+K3VypEBwB5He2MIX0TGAWp+aR8VreoeXJiteEAY4PqZ1o394zBNUaM7ouGL3ZXzxOBjt5mx/P
LZb8Y1vaw38Eu3XvCsQ/fgibMgblyOduqLs1lAS+VaNRUenDuDyDN8NnYpyXS5fm0MfZ+HqU7Th0
uTiCjISSBTACbpxELJbXfwpfRIz6qMfBCOIpmSUgdurSCx/ptb59FoG3iDZJmX3yTC/4a32VlMUf
B7UHzhJ31hSFZ6SZh0++PrpT+phmy3ZHSo+46D/BvfpjUyCowVWk9mQUunwN0AVChdT7PipZJtw+
v6T8SPNUfHc5iLcxRZJYxLYuK1Do8rtOsHPouSnS8N1H/XxBc1HtVGdlDkMZcZBIKQPxTeJ1elV6
Th0jNAGk9fJss3xgYRNRZnugbmXnhTm1vCNx30Ms71x3Zn58R0ChBTg7t4v00kOQQbxGa2wiqrIL
33zXBOIhJax/M31ILKCUnjRlRDmAFMD83MOr/47TimzwO6c9hsXX7Fa6QwWXtnl8wzDHy+GFuIZA
kGTZPlKwmUJppEoDOnwaogExKiDL1/zpoF9GnXCU198lP5PiQlu9F1SH/9pZJ3xhdXDs7DDhAoVX
12ko2BjHX3D5RVEc2RjnFin9KkibmayuxpN5M7zSHbKoW4/CeTg/1G0db6MUk8kKODVTGnXBoP+l
I6C4DxED6rupASpqt1wmvWTsWAjvoj123oHObfLMRy78i0aAjcpT5lBQzt17TwQyv7GtT4o7Lvmf
CFKDTZ0RdbCZ9E0dwl+eFzD1GaX1bfJpQd2Ym586dsxG49vex1RuI+3/P7HdG1/qvnSz+7No3IL4
i7rJ1d0dzpwqOjgFNlv+ZWQKEHoQRSJwu6jnl9ova8uydsPPqzjzOMP9SJUO8jcGhByQDYbu22GE
9Oih2juutpVlw7XOaya+fatbOetkIt2A4GXDJAZx6yOtQXzkZPfs4XPOGhBD74SIfkQMnRDyRkub
LmtYFZQDJxFFAKzOdtW++SpgqYIzLJWOnnxYQqizgRlqb4u/kZBhNmfF4ozCSaNMI25WZxP2oO50
A2ug8i7HwwvPtgIoe7kyBIJI0jAHEc5m49ZF2AyPu2vL5bv824xWrwt6k9OQb5nerxOE1XOZpcuq
4JlPKIgnPN2ERSrebFCmgASAK7RjKD8IWno2XIBxiXg3/V9kdIzGxOsz3OYr0f4UFpINTRIRKDlS
drNdJ5iVw0SrJzbdGk7cWhQdfI/poG4UTg1RdFS1TjaVG4PWaV758679De92EZzzR+Z2C14qydv5
Gs7CfUxPk38Y+Ycc4fWx1UIL3+jQRj+RntlXQV8NXlmiZZO+1xfypxxSiI94NrcVRplR62z2UAjm
dX8p+ou12I3x1aSHR9vVRyNlXbzBu0FlshUnZ4DMYasTM4x4LlAO67vGSl+DlvM77WFLztU2B+CE
7Klx9lXURrYnL7O+kCB8QaA5oSF21Lb36qf8EUoQd/fZ+vPHkJjIxgx+9AX/duisDDpf607uCgAO
/ATm9xhlWvQdyI/8EgK7livCztLq7A2NNvJPiSeQ640Ry6L7/m6rXYerZkDB4QzUjU6PL1lbvJLy
dk3eg3dKnu2q5Sryizrp5G4BwsIKnI+a8oUkdbtb20FmMZ0FinNfIJqC9CJG0a/geST3Prayzs9O
wM/s0jl4LXPsMedqlZKxnk3gtf7GUMKGHmu5su1h54uikJWECYgyU8CAv7fCUiYDD6TSdOyb5Yn6
Aqraz0NzCwz8z0uCqAynJtpd0zeHJqkyoLH6E93bMzvIJLPi5GttCuL+bSltxxlp97kbWQKuOouL
QaTzCH+kFC3VQar8GrG0FBJcfeNRiHXSXlbC9kQsXr6qzgjTgFr60vpedeHlGs659JrWdtjvwOSp
qH86oMHjFYV+Vu7BCJ0IXZL3WLDCkeDsLz4mNxEbSwTyFtu5n2Hviqk8jO9DeMtJMkZyGQXx1rBl
8owx61E0w0h8l/6C4V9OQ4QgAvNaZYE0KUhv//0LNS8oXMt22kRqkrTmWInArdJl194lUQ+CfzPi
c2alzvoAvwUWAdS3X5BkUjGhRnJ6e3kWLPNTSAVxhw+8qxSioXY71zftQ5awCDoAzKH4/lNJNpo7
7poON67/Zz+I+agVm89l78uvH4PWJcq2xnYTJaXMqI/EG8y9QcQffabdfrBrAL0CkPBp30rz8E0g
My/2403i0MwFuQ63Z+EP51Nrmh21bisWhYjm0UHNua/ZnQy7fgoCsaLw7pc6EnNJ6rwViFsw4nxo
RE2YdGjz+s517zmZOoS3iBI7oXbNKbfTaABngUXH3l3W7jLufDVIofUsilLZcDtKThgPizhl6YHL
M0VsjAPYWymDk44oUadxTkGcNO5P2pqBHTNA36JHTSavrv/bOSoL6nAFbz8mEexuM6xCDY9Zl468
6l/yDlIBbvoiSFkunfqGY8KwRcEGN4YZ0Ss5x/pc3aoH4zHchFqHNb7S3qpmsHcqoHl7LHF4tIuh
0WBueFS/+71JOphcJcgm4QEqPYk+5fHbZWv5Y6c4RWCVPwpH2alKFutMUBAJ1ou7HXyM60//cF+H
Vb19UuYcj6Q/7J3ckLj7LQGvTAtR6IUj1w5Xtq4fNC+014LyIT+BK8pxSKyFaapCMFTiF4TUd5fA
0NVphhdUhvlegPEbgF281jsGK+mwRrmpYdge/8i+R7fkFrgAclErkJ0GDNPJ7VLd2V5ax/FNhH09
G7T+Qm43E6lcWbayPdVbsfNHNNR+GqMDFrpkptAeXbxI5XRTbpT58G1Wv7zShpKSgJvFwxcYOCxz
NDBjq3oq5v07wRqF/d0NwCoaQbSC+0tWlVD6NA/irmA5+U8GJ/TzP0Ieo8sxZDaCU1uL4SJ2RDmc
3Ad3ejrmJ8uWouQF3VR9pjLcvEytSWm0HesZsuf27qV9gj8ONSzpJULoKFrH2HvNo87G/TNq8L4L
r0hGcmGmlWl4q9OiYLotYqjK3USU6MclHSTb3qbgtWwVKjkvZobiY33fLR8O4YzTvZdDP0h8MxUX
Eb8A/xnGoUR1vX23qw6/ZsEXk8dfo1VvSoQjKPDOb9sk+W+Q0Yeot3plnFb3IRNSDnFdV99Sgwc3
B3LkxoPNSq1lElIb2vlpMkajtgmYo92P0OoxG/yf87cwP3KGkFhhITWmiYYDumqnYJA7oclpYo3a
v1ByfcL1jELtQJC/5V7IGmd9caDInYYvMcJ0+fSNZNZIc6AI+HY0g2/iCxWSCq88cLkR9qdBg+x2
LyzKdLEWNw6eYqViZkoa3qefIsiYjk85TWsikyYelfCNgB6VJU0y72SqlRjFnq8uaouJK5fj1GYX
uQWIuCbvcxSMIKAbiZaJHdWqJbzvrLjSsJ9tMmDDPn7DVmd2nfmCPnSUFhmbTyIRlpJXzs6WbjkG
ztEFYCLzjn5z0SfZxGSDBdhhLARk3yKYOJPH0NY6QS5XQfOwHMvXNS0puK4btp2ss8ONnbKeJZGv
6/SguAlVzqDJ19zJeG7uhpsT4Wcp1Bd9sbDojvoOU/FzwJLMkeEZfixBuPo9VEbbdYLTUuHwo3Zc
zDabndjmjAuiQtGpLxyGuQliwfsFeXYVIF2HIHuB7H7lJAu8s8r95xEGHAfbVZscr3nMUuEVVOaK
ZrnU1vwMlpNApOLqPbZt/n1P+DGoBnudqlR3laSP4VQO1Hd5bMbXniUT6SZiQI7KtzOG51k9Dont
wkFN8RoTB8JUjey9mH/NrhAsGR67BChPzPPgOqCgDWMg4XNsfj3ZrefrW4JLiMpkdrYj5h5lNkAJ
w1t97behOVnNRc9irdSi3roJr0oJb/Z/wBoRRbA38OTSNFFkE+29gD8CJcLBbOYsVWWAS4ozf3Qs
/7a+FJZgM+E9FukatKa8hVhr9BgO+Ra9jVgzxaOtLX/i2ojQs/eLx87Mwb/F7idPIgvq+1rFSxft
qYZko4xY88vM+oTriZdg+yohCwzbfBpaySYNhK22YOyAety1M5owat3qrVMNRF11GFIZJrNQnDjO
QhKxdyTmXmzL3x6d6JQuwad7yNp2q52e0q7pd/VflL18Lcba6htnrDCld3Gmbm3OQm9LXFGzafHc
tD2VnuSJTMypUDORtkuuEj8cxy7NNoeRJUR8U255FwzSRGzb67BDzVmBSSx18KGXqdqQlOC6Ux4g
4Me5Et+SDJNZb2VaJQXOusN+IG+zNiDalWG46KzSLCCUHJx9F6rPD6bCRQZ4IoROYVJvksGN7DMd
m0E2X2PUY0ZWsWgT7rreuSYyh1aV2OfeydeojQZIuSQm5ADVze1vitpJA2XFQ5xEttAZvtmRXxtc
AfgViyjbumTSwPij7AOvl/bF9ACxFg7qlGMIytDk2+Z0MMhI9nSQ7s8z5FM75B1UoTlM0jVf75xP
ecg/Qm/clj1DVmBZm13sR1ID+lWPuGsVmyMMgvQ51u7U9r/ys67FyQxNGnrSb51FQ+rojWNZDWST
UagH4i93gJ8BKr5NXhMbaj4tVfODrG3rFVRTMpWcrsdpt0ttjtoVdAeLgGIYsruIG+LQZFDRQ7Ze
366BsxDLlqMscLhhcpUo07WhhVWzI1OLkTyhTaqpr8Spu8AXNG/z1dtcM2qYuMqvwIxOqnIa/x0a
F+T7COSXy6HDn6Ad7ZXuQZmdn044PfoTs9JZRMim+eGC20dZRv6xHclkO6XBVVydxXvfzMuO4c1F
M0ZM1kq3oVJwrdySB4E2b5gtXKetSBHcGZ9SnAMZQ4CV81NRkNhDt+kbQek5s3MTFtAMVOqbuPgY
EG0vwnBkod/xKqlNlEl/gYUXAw6Nu+8MXL0j2t+/K0nOW8zPL+SPCDOppXHZ4XfDwmK6cf5OJBeW
H+OSIUTbZcaIF7ONiZO6+Stdldtr1J6EQ5LXnbpQ04Hh+iEwQ4JpdOKbDuTi02IT2TmcaC2CgOwZ
ONveeWu09BxpQy9TrzFeSYcPoco/yGkx8oKnsKYMjXeZkVCBvq8IuhygswMYhF0F0LzoHzNQkjAu
TBA8nJK5oe/dy5QTSYZQWTC+0713KR5CRROfM3Y9VdyoUttdKCJalR7WBa7gMbhyckFZ7acS6G5z
cAwz2pVCxOtcHE+t8o8Na4jPe4QhY9VfTglb2vjXhnLkiginI0XyiR0mWpUyfad/nfMJvOIWLVc/
IxqGTvaLMGa0uC5gAFRKfscldt+kQlTFeZHg3EoPd0O9Bfy5tWTxMS4/j85BCm797fbxZN0A2gxN
4xIdhoA7YfiIOk/7NcjuhJb+iJq9ddssyiZzPp9iDhvvNtTb9IKkKQIf5y0e88UFxGZI1zc1ripH
F1pd0+ZdgOD6rBKKPiHOlv46i2TZPLjKcoKyAMxsd0RD+/seqZdPwCN64ztM3bLVr0Q8wfaZBPID
R+HP7Dxumnf5SzYS4UGAmjUx5y5ps4whp2UupvCxAkaUHgHxA3SvvsxfODUec7hERQ7fERwRoMmz
O4wTWw7p2ZJqhumhRieTPpdI3VyZWhCsF7VBhfFEzfSiU1lsYhh6h09dmYxnlENPw10I2V7+Cmf8
fTjAnDEKKZf4OcRS5usDNEp9ZeLDNpSKBXfS062be30Lag6jMFMt+7fpe2PBJCXi26WDNDr5XDi8
woxUQR2Nog+McmJosES67i8B6Sygsbz0HZfLZSF7DS/HLXEZylB6CeX0yy0L1GNDba55402jA112
78LPsETlOqdrXgc6TEUQFgrbxDEcH1AdiZ69vPqiKtTm1z3eI83v2XLds2TszOjsuA4GhlRE5gG0
eGlDJu7X1UIM8Obq4pJH2vOx1JmsmNFmRbxmb+X3uT32W6ss/v0tO/bEwo71CzdHYRZxq9N0qjDv
SueKZmbe3txkCLY4YZel+re/tfxlhjoLtXvXCQHWcjaxkGOU0kR3rN4ydAsC7R/DH5I76XlcAKP4
ynbxUJi2pjbgA77NhMGmZHqKVdDJNkoYVneVyZLfjgTPuE4t/1b+pae3fhHMKLaGGMd9nIvJnK3M
nEfooqkRdjWX3Et5NyfH8kerpx7T6YlL1i356JQfZL1JvHiXGdJpRMZaR0MB3AgZtBU2zMCPVB4y
DbgWb0dpHXBVgP0TGMGlX0EQ93agViTSAiBqV7Rd0cFENppLyoQC66LWNC7Hu+l7itDhwEskdTru
8w+Sdv4yUb9E8aFX76Whvo2HALSbBBiZ+lExIJ4jC2Y2F7UyTzMUcIPtXgKEwJdXptQ5Lxak5wWH
B2NYR28WHxCAoedEFrITzFwVdsnqxNOaClLbJ9kWjDBw7vTrAt6EBQWA/AfHXAEFL4/eNaAvw57d
3rYX17Of67aU8INIJY+MYh/v0KDQ3adhb7883ylXfLRSHZ3hcqF6rWH2MJ2fO1V1s6ZNjwz4NSp4
rUxk5NQUD6WgkLZKye7Fjr/LWjBmfXB5pSXJ4qQ3fFbNOuTP0+Y724j3lWmbuU/nWgPArqpeq5BY
U0J9LutssUKF5FN1UU434bkS2p8gfVz6vZszhgtcWfvnuXf75tiDfHSBqrKGv7q+ji8Rz5E/5PSP
xTGtVet8br6vLkaJ+XGtuMXg2EsVrFFQsHZ8TpVXqHeT2b4Y6nisNSQGvnfQlYptVCqvpDXFyuWQ
NgumQULZr8hcLdXhLCtMMsUfhJ/JBa4BpSCmA+iKJtsU+L0tVJVPsgjfFI6xQ7WuW5+y+2VQGnFQ
trsd2RDQUQ9tmJOoLyEpT+CEesrBHksFJr2rGBCLAYX4IpTBDJsNNYOxzaKUfbIVTlzwrfzxbJtf
cgy8dTDG8O08Jkt6JMIk2+D9oG1bsrhvnrPEApyQNP60ioh5ASIAb0wWHmaqf3z87gS2hHulpB25
6L7XrmJBKquQvnVf5wkQ9gfGzJt/gBqXktPtKagoW+AjZUyMvmDlLoSaym2fm/FMFWoNF6TruPbS
WARznJsJKTuEyv2M7qaRP/7Gf03DsB55NhYlxxJSE+wSj1qHb84vUKi1yK4KsZKmwsmBvMC1RQ1k
Zsv/oAY/BGj+K6dsapsdfNfadACfyW6d2Zd686WJjEMWN2c4dpiFv75CM79KIcoPA2KjFt2tpVS5
ycGQillyclhv9OVriuKPMDqsMuF6yb8Xs6i/67VVMQcPHk/6hkLApQU9mDzir1nhiTSgGgMmQ5wz
8T2Zr8alAyHw0k0ZbHILlRIz6YDvEQaX5iX5twvF5Y4hyMNMK00k9IFx3Ra7nJlGVSi1VnQTFyhW
7bk6Qdp0jNRg11X/w9iOz3FsFj+2y9PKbYPpFSChN0nKyAMWNXI0F3sPzW7N2KDQjnW/Fme9WsZ8
jU9gMSVkyLgi77mcqGzPqYapP8Hvcy5NMv8tpVKEr+BFbiOCg8LbNt5B36w6Q20pP0tBpbQEayXP
PoTzj13X/TCQv3RcAXInicp0K0qIy4Vx9tKuLUY3sH7q3QR2PYjFDg7JWtJn8lFsXws1VBoIXwXX
dfCGBWSBU2u1j+9htLfirmDtM2ONflJQHn6P+MiGQBNubV0+8xJTivVIK/PVbLg039gNkoR7793r
8SezRuNu0w8TBxlEDSfhdqKkAdLDQCAGfhbTL3Zb+3KGdjYq2W0QBPVIBBciej3HM5QJwQISkmYk
IQVWcs8WI/z9paaSWlGWYcO5D1FTsTWqFLrJLQYXnABp2XIJBD8SL6nMnhlvv71FB0GbYsaa/G0w
pFR64vSKQdqw/N8gDIRAZQz3tVmS2212kp/gt6DGAVDPDLaQipSInwfF5tnCd9j8huDFLt0/DoD0
NsZoH8Nz7CqI25Daqo6GcCEOJm6zYdP+bVY5fy0soxl1FCEKW+Kn5HUTae/qJveWvjVKazqBwzYA
mWP62mtheBn8fZKb0UhdwfgwKAYMhzocaLn216Uy0qx+/7cwINia6QZ5LYOyNmkc4GLc6PPQqSX4
Mxp2f2Ix8EnbZnkYbOT2vhms2bMiz6msolMtpUJACcjuLnpEB4weR3H+Uvnlvf9V7DyqJLG+E2Ym
iBC+Ww1sH4Kh+An+8t7CqtiUTXQcfHexcj5NUHLkK40pZgRG+8q3IUOXE4H+189fS7hmtmfllOe5
czF9Uk906TitoMJN/hWfNxSpzrooi2ndLkKeA746fVhmbPb/bolXhSlyZgoik3cAxaiB4LU02PDT
nFTeS4v+Z3RbRzQZD7Hl/3IEkgkbu7/FDfPhXJRsaZyIh9Zs3qaYhzPtjXBb34yE5sObFG18h5Z2
/vHGGNfxBP8GWaw2W1duat4ob8TtLjxCyaLm+DR2KRyL/ISt4ss7KoPDG2HPBvZwpFMtjV5MO7I6
5HC4Cxio1G3EwTJgcykkqKSPJgoWBFSjiVBNk3uaZcx2LKpye2MM9ssxL6K7mdmJIkDjI9lJT7zA
W7JkMmOEXMw8dwSyAaVOizWUE5NWhfrqYKBtOVeQe3+cuqnCCkuDph3mOzNuBbYcZoOD3cptPNIG
T9ZwHDGrIT9FeL7Ip9PVdj+MW/IpbrdcqBIx7UoBVv1xOGzZpn9XD8AEavU8JZdVFdSvMe6/bRCZ
nU51+ssQSgde+W0jvmcZf4L929s36gTjR3vtJExTIOE47yHDnjgvmNehTuWkxAYGn/LMV4tcEU9E
1z7OE3yhi7oyNS2jaajHYIU8/bU0jLnGao1DJa3rKmW71xUHRiMF4skbUvgGTClIWREtwVc17rzj
uYo12EZWu+8leLNv0ksw9BQwU39hJjp2Ou4+I1qDHq6U5Bu2liAlSRtFqtpe0ez0lhwbHk78TLhA
YqZYrQV0Q497DKBRJ4FDJEuv5SLAaPUmaR38RLk21ZJEBsw9tJv3n+yFqJ2VyNh0Fjx7qg6qBdlX
uyMNQhikk4nnfAbZj2gSEmRaPtLEaVGnoGtGURzosUhPWs4a5SQo85lC1036upC9hPndySZHB5CW
MkuNYRc0054kQmwlKzpSJRTXs/4jWUu06xEmCXvVMiPJ0kf93HxepijY04sKeArt9eSytdDGYgLw
6cGPrBDVT8bopPnXIjfViT6xFOdgpS/a2HWv35k2/9UcxXRdxcL5DSRgtiyQh1E3ULqoZ++2AxUF
F3zslym18tRIZQpDY+0UXF3nPRY90RedvNPJUfvNJjLGlFtQpHRpkfsn6sMOS/nqPn+VGDZHX7Bm
CbKtf+oZgj2DvEKhLK0PxOTTJlXATIeGX29hxJoFXREtit4fYcgcWjOVOoR/Vy/qxxtyjhMeSmTZ
3LRwlF0aqI5X3AcRTYQYnjjpsotX6i/WlQ4vISz9hjRwCsqODPc8w6Kds3jT4wqiyICdfB0OQXdQ
2TZNP9LtbaMare9SDqLYtBSdrVw+X/kH6cYjqjDCWmMDhyhmsKKPzZN3JyxgSPY0Y5czxcl2UckO
u6sLNk/pBgJAz75H9MMVikqqfIfMXnbIkPxsv+R3m9WIYa2oZ2mARfr5UD03z7c2e7tJNf5xYhBG
jJqjauEc44UzeXSuvRgYBjnGju9qwqZZQxLC0e2OAzlCbE6WBD8p4AdZcuM4kPXb9YmwBYOLLrPH
gYfv2RCbN50swKeXjeJM6hVVGIYpmtYKac8e/VfVwzyPru6voGGGjFXuwQ0Ys01sx28lCVSb9shf
CB1R4CUZ/d3a50s79xvxZJ9UEZJrD8c7oxfU/NuPdqyO7WZ8dZEh3Gzh3QkzgtLT2lpGNSjDECOt
014PZjfz+2z+aQFAWES042J7pjrZaA3iLKefvmwzid8UIIJnPD4INLrYQQOQWeF4hQo1Tg6Y9oVg
9gqnXH0SiN0xpxKj62RXv+uZRvHMbhOJV7YBwCOUuCHFE14OLNHlHorn1PkPMGYUQfpldnUAgg/Q
H0QbSLr3uX8oNLPzrctjy+UVLtKbN/B62SHLqz9vtJQBt97xneGwaKFw+jO68e7m3hyWDCrqAtMd
AnDZWmiAvKddp+UMtJvNucYcpk55Rk85CsPJC6zwq8j4arVjymvRPZGmNySmDtZyP18H5cvHTURy
k59pKaw5ePbMpWfSBVmooqS3lwvP9iEqeEdlVzMlUMoK0lfgsV98ZuMWd9M1C2odY5kcjc2PPOnm
Klofycp8EvpZ4HUptDprMRUjKP9YqolNOIltDcP+tmoo5dMzdvvkuVIRuyKNEuIk7oxaQ4Tn45bD
pQan8JQV6eOolKx9T1q2b1rAAN1tz4xRqrTPr4lxCA7no7b63ExQK/bJhSXHBnhLFxHqSqGX+rNq
ne25fm90buTSpA9DsozazZ7bRRw+9QmQOcw8UXE9WVs33tuLwpgY6n81kqcvcgvJ1gW7Kg1vFol5
IXxyjYGZLkF0/UFNmzCA4gaCZO+Kw9S78rh10Jq1MitbXKgsg2MejdkCkhcgWQTaaCPafh3mTE9W
T6cbBRTfSaToFQvNArYRrGc8g08agMC6VUm+TN2WXUZWq+RuxBwe7hBQTiQGYXV8TJcJXNYK2aaa
53F0DmKCusCo+cRDBzkGxldILA8n/VjVmaoShOn3x+osNGtehjbQ2Qrvywrf1Sn4JTv6jewgSAU8
jD/vfd5FFXYy9SQ7KqYBFhdjW/zRMxXkzFXyUUsRSp9xazr2YSVSpQMjw/QeIxDw8eHd95BPmhHO
OcH09bdVRP80AUbLGJeqSaV1nO6ASzxA+VyAwFxhffcJSKeGHQvGdrul+yUAyKJRW74D2uvqzRtC
1xgCvNVMTNXp+umRwtlgeVGIBb12iRTKiurUI3ucsEb9dHaxArn6LhHz3bX3MnxKcVT0i6FAfaeT
IC0JW1lhqdNzucJraihzZ1YSX9X4PvMbTjuCimtqC+PH9ONChhgHn8vQDcqorqjARFbx1w48bRQY
atS8lZNf5T3Nwb6yX8uc6s9Wi6pCTdW0uvb66WeP8dtqtHNsu7J2JP2G3rBDAylZCi5RgvQbSREs
TNq62OX/7FuEAZMMZYy1Nuyf0JrD/vHiVH6SbVGgJZg3uqsTGTt/xj74lCcKeRGGMwF//a/MHPGj
7BCg+JU/SRjTUWrhhXV+Wt+JIQKmBbfaitveOIFmwuI1aPQ6DYp3iulYnOK1G4rcYelxOGZRdO3Q
7pAXe/OokzhgXtnIexx+Klqfh1PIDvXhBfy7ccbTfE3XYvgOhGhp+zKsfR3VqsAPMtxLtNrmHgQC
yMo2pG2ThfrfdHsGlEdy/CB6i03GjgWqj+XOCjcYXtPrB2SJ6wJwkYY+ndNzPvfOdr6jYdFlXW42
HKJXloyAGNtbwJkUx9manZBSFi5FXJ/EqqoGAh51XPC/owZtB3VdNf/ZVflg/jLEOoS+3j8mHCa2
AGA1lGbiQ3TkhBYaKXk+zEl3pef2ZUlUJhKtKpwJJMeAq3d7dqg7m+c6ZImYLIbGzm0dJEzk2jn/
g4lRFzabguvmRVaQD2ifGcYmzDWvVM49ed44LefDRxNUCG+UxEaTQOcI5GptmiVS1n1fLnpIaYmq
4VN3aswnmgsBZBxGCGWc9qNakievjJn3gwFGE0TOoZ4z9t6uioB6N8EdoWmKKIcNGLosP/KX/OtZ
suVnDIGtrEo0Jp3rzYTabsK+0uxcZCsmtHdgwLjmTF2FwGBZX8Olp50dxY1arJ16BOJyZgq1Avqy
IY9TUgIkTDgAPTDffV2Bdh2S+KUkciJnujge7xfUMZEbGrIYMHiEzD3IqThWRRxfUAoNq8828NkU
NZOdKAmIGkCHQOatvJFdpDJJoXqeeIguM/3aYLET2Nx8cCbY7ZSYLxgQGF6gRHzv+KoyKBewBGlr
NfAtekRzl3/FQAI8F7uLLo5jujSx9U4yIAobSc47XAnlMJwz0NTB9I17mAGTiN+GVN6P+/zoP797
CdT6kuXn85DHDEuLwfU0vD0M6MKHzf21NHz7l5VFUxs3yIQsmGFnhuCunneUHH7ZVa8U8nLYo25D
V5+HvexkZI4eIjbh/gfk8pzRV7XcQF2YYYmFScg4X26/8NQIiPKA8iFyR/BmeGE8DtmpwjuPqgpM
4U8tqXZ+JkNqFEVs//ZJlEzKDfmd0llzveZoXrRoZuR19vI1onKCn5V/dCJTT3SfFKiEdTfDJN7P
b72et/b44Y8/pKZW0qYgNYveSAWypMbGtN5XTNFDbmulPVl5/quH+6TtE4iaFTFY0Annne4v+iKO
OXhEsYp66Thk1CqkabMQAfz0GfugX2RktMB+KgmT3v8Tfhpo5bbQuXQhaF5po85zijglMzirPBv4
bapdxXsUWAFlWDSqziNk6zoV0dkHc+QObJkczCIP3wQEZCiTTW8gmaj8oGvWpalo4SGMTsqsCY8X
EnewM4OKwauYXRKzrmuiu6pjgcwAAnIIqWlOvlwnzvcKwCy0/Gdv5b9fqrz+aPvycaF9RdSiy0AV
xw6dtPqmLaBq6p2hjrkwq6RW0U3k32K6VzoHrIFOQWE4TAqJE0wIpsJe9QajWQeVZ01+7oyULpEb
9g+z4+cMExdLhpERtVOQKmCUE6YDXpLT9/0AfU5A+p18kb/gkmnUFQzRH8nPIc1UsxvwsU9Qvb7X
1QJkRhAlBaNgb4h4i/ozpyX5NxdxhLw4X7Rua2ufK8QfO7JScf3zhTlEud011lLYL2+xamw0h/lW
o1138IQ4AUgMgBUOifvfhoqVa0G7hMBiOLJ/yFkVDMjy3xpQ4Tn1cLk3+eFfAfetOWX7esg7f8wY
w+wftKokHGSoX/P0HDW4anHRxXJ3neay1nsrzQTFqXZZrczIz0B+riEY1oF5rhIjufJ5rtqz1Fpz
T5VQJXey/M7sHdFB+8NjXcCZ7m/wdxyLLHra+lqUPvlGmVLADzqH287FhRTVVrG/vXoH/cze/Zr8
rvvDKlV1cDG5VlD2hmrR82owIz6Am7TV60BHzPL8RXxIE6xcKgAigEiJNQLNlApPYXQMi514K/1L
+URRJMSKa9vaJUII6Yd+9y86gV2XhzqrLwD8WURiFWGyICJupa13GGC1beXcFs6vSWRIuRmEJ883
+QMBvLGOa3qE0CI7NHOYUfGKWKxvqp7sGFYgaU0fFwG9paY+MhEBe3rQzgTMgqnvriBrclTzxFXT
5uurSzMRryeqFdpXqieezYjSQg0xD3rM61KtusqQnoA3X7n1Jx05JrLtk0FpjIJIs/ApaiHozlyF
r3kBcjTnp6ZVvioYgFPpGh2ZHK76DiM3CZH0a/F89AJou02dpMlCrUPcr/GHxpoQ1/X5pSvCoBEA
nCozzktGQw68pHD1RilFQmIN4Yi/xugcjqepRCKCxpqX4P5Jo+qVE3nmlWrmUaT8ehba+rxVrJGp
JbkZ5Pr/Wra4MWG5hLVe76BC+P0a3Q1QAcd4UTC/pYubfNzMfBtkgK9k7YHOLmT0gVXiM05qnx9F
FchZLXFscMITmrCt8gTTmu46SXx9USoa/wU794S//+bvipg7H6OUgwopXRcq9yIhEB0kuoZxbS1X
rFer9obeQkDcckX0P+KnMcJ6SVZB2RqHG+oOho1mJoQHBVFaP0+h1fkp3nPBypPo3QCaQ034VgJI
b5Mlyw2EgA7VI5/+ek5PyVv0l7lGCzvCKOMejFZBZxR7gt8cJJ+GblwoVPee0+gHc9p+L7hXu/E0
WNF2KhQ81vAs4nYMMzLi08tNNkjE59Yg/Nm3IoCs1twOOj51lJdvUQPExwgLJ+sk/a92Vm1xIHfe
GCvyy1ZfAh0PJ6soN8gU/dwtQwg6SUSCSneS9bAgneeVV3PRPXXWBxrHERbNfO3fKeU3lcsJ9HVz
VerLs1K5u9ssJGxPt1Zm4x6U5m1jeeWQOU38Sd0Xr9XVrIP9tMlgsuYhnubb3alwl8+XotMi8UW3
PYhUhoEq7bEqEa9VM4zF0SOX6JCFD/o3kyDonTXEJhcRawh8BJwiLWQFoezedZxYLa32ce0eaxkg
UZ3tRhnV1UQN8JgTTEuWi4M011HKrqurWDxopZTFaXAj2faE96/2STKDzhi3uro5Tx209f8BjkGs
uz3vr655alTOd+VrwSo2vvRp76+TMihtvzd3EwSkgXFBuRwJdeVd38wgdUxPuVz1VPmbKf7kNnIc
qoI4Xxya9uFId7AD8YXDkf3VPioQNc7bv6hLy7PJez7BRuZBzfDPNF29Lj4pd8vD5eNdra9YAly6
02hYXdSua6iIlvyEWPKTXIT0FMSWWbxN74+9MHMrhw6tBnLf3ftL0GD6GLtHZ8xbLz+6HWMcGqLR
cZjOS1sh2BOfFuFIriVvx7e5E4JqHgUu3+ORGHJ+FEqD/uI3afkiA3ft6I2NqVpxq8fwAnDLCo4M
1ch+0rmz03P5fMGtu5LhYDEMyPJGiN0YksC2psgXqb7Yu3+WvzrI/Te3wlPskO2gVrjHkAPvXCmo
3zYenFxwFBajXoY8Y3oL6y59kfvu9rN8sHfOm5rkwLKrJOAUrVoPs0rX9Otg2ZED8z0phYMZWSxE
nFwZgaISH31OBBl3lFCCayyx30ddm51ZlQr3OBE7RlqQ1jaV426uearuoa91HJtudsqzpxCukrh9
14CcHRfsNhuLF356qWeLfTSP+KfMS/wC7ELKAih5HcL0WS2vwqEK7e5v5xL7y9sLhpnFXOio6Way
+Qd1+v1qNfPXd/Jn1e/yZdcsCwx+qoSuVqlZFTPtaxznP3sU7lTjWysbYGIsB5E6uc2wumoUAvJN
GXcAXS1HgPM+ZalngbeMbMBi3UupCGqG4MHFM96riNdNP3UrEDsrRZoqmzqyDQkiGaWIlqV6ucKA
5veTrgvN9IleexMDX1cQtXyOGe0VP62w8JRE/VmCb8UpSn37K4p6/jTsARK3dMWa11zO4YJcRc7Y
Wex9CMgGQw3Pqe5gDDT2mL2VOeBT8BGNd2oMQdcifFguEFTzh6tzgPjaMsgAf7b5PIrLVwMFignk
DNS0lk4y0lrVh6qMnwbjMpG54HNPbyGmFZx7HS//N8POg0XM1iEXqAHsKKKQYzO7ld41qH0CriO4
a/CBb0gm8nkoNPsXTw/SjDdpx6myUoC9xwmETXeVr50evq+uuWfSOp2EHgOb1ItmDf499uit93MH
5+b5CeHLSDmbURVYHQ5/7Y9aTNeTC049BfaCKJ/FdRhrgIavathtPkM8Nm1GswHIFb8WdbHaS6U/
9MrnNK+jYBsYCpfECX0zBa6famOAcLKsH9yjuEul//MU170f+EDM4DrsYHmd1J5DHG0hWbWZgjQf
XgZ7RfVgR1HEIVC4CwYOvO3YFRCUG2YQWl2YxZWtC+rh8K4LOTP8kaF62FQugXR4Ud60fq9gmAlk
HytOfxpwoKYtnxi2uRZ/l1YgUmVI4s+RYlARg6aNOohqNejNQEYzrxTFp3aqyLVUt1uHOYlKR9nA
mSB7prbZeY5n91LCUsaVQTBSTSFFUHcQsWb4SiIZ7EBFaL9czKX1T1aXgT+1vYqY/O+LVt/WF0N4
pX48k3kAcyQR74Nu1YJcOB47LExwsS8KIukraqf3mJW9979Y7swE8LLW/gOQ7e+h6BcdzRYwVNff
OmZ5Rak27Kq3cRTZhRiMe4jlk/8rjULFPH4AUgLbzSOKiG1liFKLJoodqhNky5ntXi+zar3vSoz0
uIp3k+8pYHDPeqAnbLpnWDaSn0u0BpXCEdg9eNgB8OZmFePoF0qi9kCSvo9xIEUNQSDsCoVZCFx9
AxJkK3w/pXq1SWDrakyNEcEj0XuoaMzsptpa0FWZ7/CJylzaiaOp2dRNykPV0HNWtXN1XmDDcg4r
YNdq6ZjdGKhZWeph7gTBe23vzCEkYL1TGCmJm+pm269UAHRr/TV6a+KMi6TB19SYoNf6tDYo9leo
LikjVNKDv23ldnXkOQ5xXc1g+/7+xbg+WNHojZHrm4HNweC3eXzVO3lwZKpGXg+xD4U956Sxifn0
zl2Fq5qCHC2c2EjozDIlJiZ1U6x2z7L76uHUDQdhHBgDLPpCbIDo2Ng/WiwwlXr5KLpNHPBD1WKB
aY/oVvbJ6KTlQk+cn5IXVJ/AElook/OhpYE5vyNmXRT3UsTnLRJUSct3HO+Nh3ibG5Ie1POO7mfX
qWrnPFSd/e7pss3Pyx1MzdVzAA7Jqjq974vSWajsAAtF7+ye15VXUQIOBTe+GfVRpRb4UsTyaS72
hMfEguWGBvJlF0kttGsrOeGJmJKvolvxFNAjeSGx4s8YWTgTilVzhhjnldXJIq/tOWHvBE9JXszl
RKwI7phPTn42+C29kUMs0CYWAlKgM2TWKQGxEdoKaF3AdQbXxEyk1D9mADHKpRZgq8SXG650kBcA
T6Sa7pkcmdXG3GW8gSBey3Ql0AqWJk0MKld5SkcazPlZj16KeQn+R0m+EXCt/5JqaA8AhJv9f9yL
EVAlV8f4LpeoXVEyzsVKCmyoXKxXcqweYxx4xS34R7fYj+Q52jT6DnSzksWisI5zS64jlqQiCoFM
IVlabCZIbINEtEh3nqPJopSpnEFNwBETlL76MCow58sPZQV3rYqgI7tYvsgC6ZnKm6hMM+hbl8L6
gZeOkiCFFftY/Bd59DkWb2yfzqiRndkNCYpGPHlurUNxX5dzRHWkDhJygrOU+Vm0L5kQpBpY38/z
qGy06BlHusb9SZCI05fbUj9BEV2SKHqIWvMuriuYOCpoFo2e5buL5VFxERAjzio1I2ddAxcP1icg
5MJWm3k6vUVCe98bzTIYhrfE/RgyRZLUPvCEx1xCEoGoboOv51AE047iboDkycZm8TVgDk+gzbFA
R/R77pyUqWDOLX8nsDF4c4+D05oCMlKONKeBHYCpIn6dBINX5VmH9BKXjgdItgNWs6dzuCWpmfRG
ad788EzBnaeolCd5XHeV9EK+GeWlaEIhQMGvKvqXApyZcZmF12TtHaLiupbt2V0EMD9zzU07wsT+
4FQLyK9UK6AhjEPceEQhRCrTc+okLDobzKoxeTyXAOtq/akmyM9rYkAgRibUL+wTmdQsz81T4GAZ
dXRcEOB9luB5v95Lsx/6i8t6CbbcPPUGNuD1xP8EnbgHf/desBxbEuYMgiO0sCMqmvT0t2IBl0za
5S9/UycG9ygQTQSBiZE8WztcHmDHPcSWKyRVc/ovduX1z01JUExNob5PAy8N42qAAeF284q+uuLL
yNcyI2PRsQobucKDEOQDqNU9tdJMeCmpWWq4sDU3MFEIOTFY66A/ybNFhBhrCROcky1k5ZMS/S1k
Yz4yzgn0XEr3BrHc4ed53si3ejJIPZKio2fZEATtSlxO1fftf8jeUgQLL9Dr6pDQYR4yfjLwhkoA
YXmfSra/19I0aQht7zi2YQ6DhLVcf3LSZWGfJmBPDyceuSwwzZclgC0yl0q+UhBavygyW4q0p5yS
qYfEYPna8eJDqOiIJYdSLipSutGdtoOyhKpsELiuIjnzZFlD9130XJfcPyWhTkgqCaKj3AydfCo0
823857j9RvjtsA4q4764jxeeAQInY8ckw/hu+n1Of5/fyArhbS8JgIZ0zqAftKpwttvnDN3QHu+G
jLjr0Q5f4c39i24U6InDOJU7roIzJOfHuErhKIflRCHudh+00fVIm4sP56ibiSN++JmmGoLlbgoF
i4axu3oq9gZ0CuXy0Q073K6I/7xjJa8G/WRcSzZUfkFQGCF79WTmM22g2Ve5YrQjhwb0/c4A4LBa
C1E1KX+FhOypZhsfi7URYdKgSMPxvVnCWvlZfccGeBR8BFd4H4gN/s2EeNUFjrcClAU95qEXNEV7
0n4wIqJ52celFkdAQrqUESiIX2IWlBfjFJvvvQz5cGDbVRi8+WRSWZOtViLhkjtuKad/moXoTksC
7nce1EGiRvxfkzOVLjpnA2hGmpuT+M6+D0WJmSm0ZEf0zHNqq0RzHlFPnOFci2sWjtn/0vYqO1UZ
yaLhERi/me4iUrMczNUzn4p/2F9HbVNhdBtT6JAyiqbajF5mjaGPbcH7RQ+ECF5iRBWChxV2W8Rx
Qo0BuHGryWTsPLYZVysjp2i/xyj1SY9Hz7IKhIQOWqNRDE77WJdpdS9FWtFFV+M3qeobo0YCnxIH
93mByuYCrRQqt0jCkBztUe3ekaVWiktVi1Md2lRoIQg0eiqRopVnOjXB32RKXpqwX13XG4JpaM3I
3UrzqlGZ7F06qvRAr+Bsxw/ZsynBcP/0xHxD6KSkWXXK9RXk6qXdKBqdBWsOlDuMosSVid3lzsuq
J1EuwYf6Z7muRlKsJQnNc9IVNQ0bDMf4K7qHqWkQOVPtW+b1f6Yf99AFCKrEZdIdLOZLU8mFcIN7
JPKq9dWvJw9WMeVpnL3PfKegKS9VAB11NS9HPIQvk6y0b8U45eHYDyvQBB1RbZvBq3SPmAGyl0f3
yMCkwNHzZfYAXAcjA0hy0VhuuSvfEJiYF6ta+Q/ZPha6UDUUzzfT4HPAHWx7jhR03WV7UStBBH0c
aCExs56DrHQuN9+t4Z2KdFz9rju0ChKf6agpplmaQgpCv2xTWMAMjExBKWVjo4BUtJb2pBN/dpQa
g5pTZ7vMWbAVmS5ipI74bufGElRekdLuKAh45BfnXEJ3MEG5KWZIrtZ8PybZ3oQT8sLXSkSgrw/l
VxDRC1Zblr6teuRtN4HMilnTRk4gTRZ0H8xWtkKIueQs2lTOhoDFx0h39n0KGsCVBCedcVeRY3nz
urWHZpjL8tuBZChwNuiKRC9nA0++OeNw0mNd1s2o2r7C0w4iprG+VE7W28StkYnBR7lwA85Vvvhw
qFfvrVv7utz5MbwFcnTPwpX0kvEM/Jy/exRQS3QLY5B3SDxkV9uLKjFgHMwXi1XflueiC1YAA/v1
xgJi4PAqKd6ZGmr9LRZcGmS0hvze4y24psjZuBUu4tENxUCmiznM4GY6fddnstmAEiIpelXOWmK4
f0jkYLypFnteHmU5gPVYGgi1wevjSl2Xv7fJN2lMGU9k8KrtLKQpEVmZkIuGPP7xEfdKRrk7X+r2
N1JxGU7CbzzO4DnmmVzgUkw4Do2gHFyFiS8eDm2X60qSwBK5kkGYDNDIjt0EgE0uTGp5I8PIOBJs
bF79IW3O9+2kTxZaPmGx0ZpEVd+Wqk/wihqGmVG3wnWTIOJxMEupMOSsHovxHVc1ipaqFd203ObH
bkhXWrrRejr60LdGvsmbyN892ZS4loEKmbc1PUngHPCOp7WrVe253ux1j3ASi6Nf2dMJ2MxwbnuN
hdIxEuY6k089Xsmu69FXG9wD5JwPypl3agBgMYLI9o7XAhCRN+KASvuWV/kyRKwGFB2rYsf6fYhD
yS0n8b6/d72n7VP6bevyGOnLVJZIbRwC6qi7x2aE+dpupGpoAsaB6xzeOeIn7++YZwsra3Eyz3zF
Imq4Qjv//kIVKgn0QRjN0JFYv9OGgnFE0Yef+mXEdoTdzI0q4qhF2uvm5Ymudc11CycM8ueljh6U
/wnysxIdelowc+8VlaeyMhncPsUmNzKFirr1Bz8kX2GgM6Cbqjs+j/WB0BgxkYaIawQm2Yy/ilkD
I8vJKsGPR732mZE6e9LHLjKQvCOxVnyYYFStQwmPCz3zZXg1q7sr6IcrgPY4KlHTZuejBU8Iw8q0
cqiEKRZjUpKJk7A4aQW/E3NmMKro1hk2NvZSFxb+ahv4GseEqpKd3Gk7N+zFUjLyzMpCBcQK8i7V
TmSaJjwMHi5QwQw7dQVD+XkUD3GUCkFhlvMhu0or6rZhIB1NjD5TrMiLuxgXb64EnrSVFHdVNpy9
RtVFm5OESax3mKt+qlFOGMCArnGGBrxIqiJ6KbIRfe+UiGkFy3WiN+PSEsc0BPjpbp8pgB/7LqG8
+5WyWLwhLWkR/xBWU6CvzGcmvA9+F1y8mF1CloNSYEbGIL8wNRbZ2TE6ycsLJAnC8XsUqYVM/g9m
Dbq55PMIlxYEExhL6l58fLruwC1TEfrhYzN2Xmuo59Jxd9n0FyCU/ujkTE25t47WSpLj8ocrNM12
kwwQ0oQi5qkUvRk26d5iei11HYwM9TSUkSOWfIERow8Lqx2kS48bMujjAW8i48bj0seItkkoYOIz
8xRJm2V0cTvRT5ETVOxHp4OZdakKAj5AXJWsv0eUjFTECuh88sP2y/Baai1gtKi4DVXXuEOsiBVU
QjoLZ+Dcegmp53PdLnl1uVuceS5NYbg48Kx3CYUl+j03P3S9sRlqZXGr7H079vKwldwdUUbiqESp
864gd9GPzHfriibUqTvOEUjzwRCRmu8pnRJ5HpP/VMKmQkEArX3w/EJ1u6Czb9nCXAYqtRifFcnC
uDhumuyzkAAyK5IgAuPX0zx5RqYOaLUskVRYOFAVYFlJCdLuRF9FlU4tmeUnKs+osWo0bHwkG3J1
Dlox+8O0Q9eV7zSIChT0J67hOHWSWHal1ZLfwqqXbVOTdZ8ffcHZqfxVzeLQqdw40076KRkMdQpn
mw4FxtCp0vHCN3dZOdCUKocYhI4/QTApW3pScKI/pDK3h3LYmT5Xau7U7sWKNr8QUPMmjN+GXo7S
35+6CQZQ3E/luyIUAiObOZe0VnmR3dy00eMB4W5T6YYy5my87y0kOklKMi8GcfJ/DxB/hZlSi9Lx
zJGEu2jw0IXsnSHckys8AcqElsOZLlBlM+OhabZ5ZKN7yVCcqiSZy6ah8K2KkYE4BMdsYb+eD2Sp
vOlBgwW71MZJm4reZLfSgIgCPfrx25C2iqm6LoqsqWDkZ/3zbXZQSgBC2Uw1UxSkHJEoe7ImvJ1X
qLsoxF0Uk/t+TRIGV3t9cBGNEtFz5945S1BCKUSsIDXAvh4pyuIR6R79+FY1E/wZHj9JFhPyES2g
P79+HMT3jfRKCCAeP9hHXN/1IBbSGS+oaOyrJGOK+u1LLx+svSnlLlSjk8olmOf96cxxqX/SIbZB
3ORv5xVumod33+iCeNJnWX01tDcai3ND8WPz5p25756zF5u4tqDagK7t0Gj0Wj52D8MKy+o6Xt96
r4tQ8Zw/EGx6HDz9CEHORnlx5iZMiBgywDSnFc0CCBiTdespnN8+4A6w4ppj8o2NM3ny1rZ6oLD8
Qoo+/GK3dXrOqInXXg/dTvI80U2xuU1rVs79kmAHUepkEobXhnBttHCDp1LlJe5l5o5eoE7UZhKh
EzKW6xjiJj+wvL4dKad1qDLM2I/e4iANwE+PxdS0WlVmJYvhDadzM8b18jFYpant99wrzH7bPieT
GIz2aUNawEPsy2l9AmLT9QCGQ3Ls5nP+vRqedMaKM7PrFYSyBNh7EdblPkDnUa7zh1YV1L5i96RF
HcuFtE8YTcHMXDQpWDTuutAPeWVD5pe9iJawLhkjojboI9cQjrdINGsVNbEQa7G6UlIJe39MHo1b
kqhe5JnbeNWwn5vBPOjQYp0V30K17R85RePwUghKlHYLuf2p62FW7Kr8xGpYDUpVJiktVMHCsGmn
5kK3dMKR6G/imKMVZX69iSaw42zr96xZRqPKNCIKN9wFvLhX0RxT4P8aXP7q9RmQt8FuHHs2H01o
sClO0yDxtnFdoy5eEKzLVfxsoJDlT5zS+xmVBwYP6oN+sKomYop3I0m4bX0WJZO1TMYFNZtR2FAT
ksuYQK+NW6zgmJfwGX3+pl+jbiFk9e+kd373OuyneAeHogVmqUkp9D0RegnMvcWbKP8/L2zXtK89
TUeFWvuNOo+8fQ30g9vzVt0k8kyl1zRkpujtxWYvi9PfoeiYxCZsdmJPrCAOMDfXEYRdJJ2Vkon5
yMKWfkRiYeAblTfjQu+b/xLBQKEMD/nVzBuecMGy2wyesVYBMtb/w47k2aMuNPmiSYj+USkQjZfF
J15MYczOEJSpJ73iMQCytziGMhn/hoHZFXm9h4VWJtb1E+O5wchddKfuNjRP9bGcccsowG7qTtx7
ttvxSDcecEjikgrmKmPCwOHVACgvl7ciwPbwVGIcBUhAYilzqdn/pxkNaam1/i1S/a7sEGqE/9BM
zJGpEMAu5q6PJXuEaUwhoBApMPYKlfjgX+bityLen8D4a8BX16lhVF5Scjb1LwSCvZwsEU5kdPxX
QAf+erdN2W+4Wd4MTVHIOANC15u0BnrDE0VweaADCiyButUuW8lKbF6hSQzN1Tn8gByGCbJ4HOoe
jcM9L4+mbvt6+F5Q9fwNJCEYXpukJ2VYn1Tbcg+4Ie9O0rcjRaLuL/HJOim8XQbrTVNJdAHKCBJY
HtvuyrSBrH4AHn1YPec+xHTVCsEmyFvru7rIfRX2CGXPhtEoFXPtOX0nwCZ+JAZt65C7YqaaKCsF
m/kO18An2xWBxFdLs1R3CK9ryBABqSHmOrVqfOk4f62fZAm3UNonAZn855T/TXdkw/4QgGcVOPBf
QAfL5O9oKScmGPLkNVeRObEGwPGy3cVaI/OwKDty8Ur9k8p51egHRLuxXWWON4603txHo70rTLrW
mqsCXAnFl1NHosjCJ+OA0YKiu/BoFR4Ql/sJrGpWZoyogVPk8ciEm5wmcQpvSE/tE7yiEn6ojgsN
VMGohKvuF5c0DcY+X3b1+EUpSo1reaLImKYym/LX9y4bWUYX3v3er7DWhUGQWYbgj3Q7HtXlc577
7DW5dWWDD0J4AmRNAlizFIu9gQ9kqo/g7+T+gvrdAQcG1TmjpyzGv8Qt+fzjkojQaEq0KqVjkOEr
W5d6DOk8beomDIsV1ngLgJf/Mjsm62i5eA5s6orwc4JT2koECGINsk22RsoCZG1udKoYpuqnGt1y
jyz2ebjGV+hzeuQvDuk9rv2PP2pSz3jAMuTY0tdY5jSxqMy0Uwu4u/yaupBMmW8UlS9qThXZiNIH
fft0qvRTTqBhR5DVLal3u7uk9iy9f/f1xD+C3Z1sepUTYBxrm+Dn7Cv81ah1BLIUvUac/x/FtRWb
tP7Y3DAD09FrUYNApzFMEbeBiH5u/Z5WSGXMdF5Cg9isooa01n/fT3GWeeeuE6AflSInZkhM2BqJ
fBVQtXefP4qz660iimGr4T2X8sETBe8TeOLL66DFvvRdd1s4KHLvwxFJFRfeznEyeeS+7s2B9CaC
YPoHAhm8Ryje9kYd+/a/1Thkmyo/3kF2ZX9dHB5KqRj5YPvQFPdEIAEPcvzVUGVp98cLJKYoRA5/
ff4Iyzay+siZSz7ZA/4Q2Lr4qpx6VscmNYAM72qp5D5pFMekNN5F3pyIRcSDC46tEIOWo5FoGtfR
Z4H+AmP6/DMBzBy7A5po1B5AXQSD25sEpWF/mM7Jdp42EOrDUj+991rshKAu/xCgjzXFHqjGRaHG
odvan+bKyIeDCj1V/0GJKiN8DDapWBkc7DsEeaKBe0LtMptJbAbh72AuODNNXuAN7hYUpZKmTD/5
sYmlWjHyeR+1zAh4MxUhE30JDwtm/cjkuP92gRe7nKiqIVyIbgwL1CZb2dLSAXHgKLsWeULgQrhT
FQmBAHjfMq4ad9CUPY7J4Y3TNTrRqy6x5w+RWhV0EImsCigDs2L9KJxo54j2K7op7h9va5XsreLb
7DcNVpMzcAO8Uaxh9KlAL4P7hh2aveA9eJ1pljPg2UBCRc2igu9cTXEhiIsquIpEfsiGW4h72xQv
WgJ3VhM+aaHgU2vIcU7DPLCrDuvfjcuNg5GYkWet16EktxKw2gPyQqiVQ5zfB4YTmNOejekpLMRC
rDvh/mkgWMioJNGX2TYIpPzt2kUfIRsOfwDq1+NFLKnKYY/8HZ2UbDWjBiOaYLrAzgqTwVvCamvn
r8VP1ZEAZfG0vwkH0xyrjT7s+id0OO0tGT7Iu6p0AB9fuS6wTmyk0A6lU86Dcw3XThEeAnyljbL7
cpAXDTcXGZ7VQPiAfK19aB8X61AWNm0izAh/3NknVgdlYzH4PdHAhtML6jnl4X75YHpjDlKJCDdU
8RgE6rkqeZe6i+RYW91o54buXAKwEWGjjO1PUHB2ro1PPB42hlYYYe94XETlh1/z0civPVny5Icv
q2unh9YUy0S1TWR12pHQk/9aZG8ap/SzoYHfr6s5x6AxCrkfXwA3TPHjONUKzKSiCzPYYpJY1lra
sP3QTn96IAZJV3xt07t6cvKWzd+pHrtKBgwnWZd1l/zsovHOI5Uy/RO7c5NOi8bFoug+nE4KIauE
Yu1FI6iEW6ZK366cwvJVWQQwafu6Tq1m3D08R7V1EW09k0EiYi/nScfkYOQB+kjinoOjWMF05m6T
/c99iipDxNc6AbQSs/qO4mFiOCY4HuoODbpIO74IcbkKTqQ3Y/Y2DxHJa5PJ56kH+qEVCETGWNrF
+yeAa/+n+NDyB/Fz/5FnqZWwqcJX/MgdpVa/mN1y6nxmRAO6ikwbZnXDQEaQuYrytmh9zL3XkVRb
YU/aQlo5P7FbbxG7x2bP/+GhduH+i8I3Rz/gWvIU39hQg7ybWCBg9XyLEJ4pCIG6VjqpmsyZQzUZ
p+uOEseYb9CqLsUTo2RTZuMoYNxmYx8+A3gwmGnCHT8rh9IoBtdSHmbg8Q4jKpHestj/dGarX+WX
rVhyhzzD1D0zb4lTAIPiz3kQpf+lvBq0doUmHDArMHQGIdIiA2PCK80hpnPiwwzxT01TZT1tZksF
FFIZ9jUSEEgoRxDoO8MYURbmSqg3peR9G1T1VVBU1uHhR2yhxahHXdT5ARlSPqN1B24DniYu1qex
4dLSgcotU4q4l+kKy7qGgadjEjV0yB50SmQm+v1Es7XxvHGhecL1BuX4udB9otMaPYQZ7RyFytJe
miII3b7WDuVQSff+OJJ3qcBBgpX3X8wv/np0RmHcwe5gYCmee+PwlYgSucyXsI2FHCVRNkjf4sfP
Ms1Zw3sALFRej/ihEhXRRtQShdlrLiZe6WJgPBYdJq8WXGHCU415XEMowhNTAaOhpDb3tfnWqV0t
1KUywlrJ0F5JJ6rVrbFl+yDprQCFJX5hNa15jUnr5Gdudkd6Kx8S/VERLNMM4AZ0YsxtmcKTZoe4
6BWys28WMk7c0/QuEs5I/Y1Gj9r9FWsMl1Fb/Df1Nn/rUQ1p+2mcqqEWtESsMT6qukeqNCb/rXOZ
XL8mTYUXTJtcT+yGATaIIP72SpPys3Uhv0Q/VyyQcZz9PaTGg/36DvbzIWFnQPvGg4w7XeP0v9Y2
z/TU4onYRdnd2kNNERI8aGkavi+bMlLrG6rQKCIOMpJ+6aPNbhdgmqGWWMhpQVlnyzc1KJLDu8/z
9MaMFDrUMxfD6yFQRnEjLfLyvPs+6KHDwVv+qNr3t7dcqlQTuGYY1ZspstB0Ib+FFGR7dtSzOgPW
HGiccCYZUTZ6Jq10Yfn5X52AWMNZ6oWMaUrz0fiLJgu108mmrPp+/B9koIT7Soelpj7dNsqe5JRI
7Z2vWRlDSvPqj/zoI35uB8kFCU4Mj/G3Md8Kk1aUpbmWvMIW0NeAbiYxaxmma4C+/Sgqx3WokuNG
9SrOjNZiavjf5Wgzwr//e3gZilGhFpKYz1TrwIgIl/bc9AbRt/C3KToIdpnr4ZJOtxWjT97kGIYU
pfZ7MOsN+jlRo/3apetBZqnmilGhFr+qxtFTAEiKUyhv2FxOvc3EREjj1a5/uMI31BHv1bBlB0g3
ZtLBo6NTON3z3BKgZ/0UDshyORui/k8M9ZmJUIY06OhzQdapHEVLSOdYcah6LjRl+KEh4/ASGf/5
m6xKjHu+h24O7b0g9af53DaxwTAfExsVmQkIvfX6Y7AKQVoq4x8jYIkzho3s7cZ/w6Oopk3G9/Fr
Jp3HlnjST27Y3LkZzbmmYPj/dnf/nYrshafOp0BnPcy4ahbBp7v7/TlaMr4QCg82XqsaCe0VnvqU
mrE5GnMOqpWJOO8X5MpMtVg3jUR2sy8XFDTjy/Z4w8I9srVVSGlECfwVYCUi5lq9HcrkzIjhoz6y
O0WrNil+MRlhREvzYgGIDiBOQFGYI3q2x8hIhe84ykQKRNz355Ddgw0c/P3ecewjTmGWGJoJo1gl
Pavw8q6hfnN5HLlQ+rcoAGjylhRGCDTkGsSO7/0o1lBGtbJAxB1NNyja+N0DVxn4L+1ofcp5eRj7
OGxy34BePw+W1OqrlpdHUkQ9bvc87+xsnbUttagx4nd07cZUT6LNyEpGCbA0k53tCfyYbWzC2M0X
IZzI9jzFdz29wKoE1pW6RjsbGSTuhdO8n2o9tEIkZFvqIUZdVLYivf5usBbgZ9+xogIvltiDboHu
mlH8TRfrAs7wy/1Tmg2m99OsUGHZctruKL9oqXRykkgNBBXI+zKQqpdNDh/Z5av7pdJ3p5bt2JnI
OXpnOBrX+MwRDn7u5/7WGn42uwp04R344dMxOrsP76VjsW8fWwp7rKx+q5+NNME959DIbQoY48XA
LUkZmRT3fvOL+FpOoeZUQL4Cxqvp+v4okxldBteJrD0nfGOuuAcTgR8ACJrhaIy56yJlXyf4I9X/
bOdfMGmz+ziZHZ/vDsLN8W1isKWqviugnFbh3Kybcv/IFQrCJHf7CFRXMKozaB1tP8EYfdLc/pvu
gdXIDriXDgtV30/b/z/aD/5s71YsWJCOaAm6RBh4xHZuERT3sKUM4PRyIlU1T/o6j8IVeK3P8DLP
tlK4hyuhl6FJv/J1r8E1bOTvnUry3952lL/mdAKS5aIsADzk5oGL1+914y/kISBlZLPsQj2x11XK
w28W+LI/Qq3zxbAOL0FxXZrB+Sx2ckxN+Ob2S/ctYaWZJlO6+nEaebdXo7jfKM/VDToa9OEHt+R/
zDsdEtJelF1gPVPoAqv8JoF22iKjzJybIduOIYTTWvO35zHW1Ml5YPv9+Qzue29H5KWwK6e7ylfS
PrF9sJ0bR/b20ZaxP9u124qeJKJBkbE0gL2G7UKJitFmQi4Lv4b9sMJlG2Da7Rkgy4eO6899Ysb+
Gf7Bi+YXVAvPXq4lEKlWQSu0qnHD7wd5F5DCVTU608yMiApKKjUlUgDVWDTwraN8XirNkb9gKo+u
hHfX566RB75UVn2FtxDzrey19YwlqeC/9B49UAJgY/1k56VWZkMGl1TV8IININkkWOZGawl9sI7I
W7GY38UjSCsrAXE4VdwiW5R1m0m9U7TBk34KaLsm5W7A+d4jj7wjlf+NGGPalsRwp4IAEIX8OUN0
dUJWwRGkJ1PVYzzAKhPtBrCWYx0jbtW5dQubf90BSs2cYuOq2VsRRh9Y0RrYHd+kxlSjxs91HNww
URRhUcj47KyikP/r2inNls2HwzvpqTz/2nl6Ib6ysE7c1wcxWPpN+ogVwOAYZ8zKGrkCfSAHWsOu
s2fVHq90810P7hnl5xVWB06XgPiEfHoKL5ygwxDB7STbIrJa1vEaRXkVlL0XIG0IlG18LTm+2LpR
2bRra9nIX1SGe2GgSGI29dfOKum/v6anm+4Cn/D39CR6V1aJH8yOfP05ETCX3oPt+KOAu+IFuRs4
Iw7oRa/isgK7tNt0Cky4ABqevhkw1DWrod3Jy6ycX1S6Pxv4zehde1VP6q+imNWbbUwsF0wdWMt7
mJambWEta0JdkXKnQwNQ7f912+9GNjJL8v0hnfTWz3DmE0k81j5V6IM6sY466yYXlwjXS3LnGG+S
bpg41+B+RamHCHnl8aYE/+lvdzsIBIQ5w0IUW4H1Y8KOthIQiZzfqAB3ITROz1T5fYp21wQn72bh
geIbvmoPkavXSTri8mSKIARaix2Ui9b8UhfYSr2rWsF9QHoXaFmEt0PtGK72WQwfczkQfUfMtRlv
kk8kHh5T+53gbCx4SON4z5/hti52Bu/78B0KmI6JUB82igi/FI7eIGK5Rf0NNSjiGW7H0irMRsjM
VabjsK81XYDAmSp6tb85UIxphm6hwsYy3tKOGNkFliSHU/BIOh+JnZdYhU/lThuMFawKHZZPsMYE
8qSJL+Q4h+w4C36LLoof5OpxmfIraMk0+7zH47QW3Dp/pWJuv3cuCClQbnlvtWoGiKdwNVfwxsbh
NXlSCxgDA3lIop/PJEHEB5x4iGb6JCpmEzIMTvobQRYzTrQXMIyJf5UGC0cFM5BP9RbRiT3rp5EI
Ei6arfkwMH9MtNNaVwIWOeFqIeVWBAe+tMyj8/JuaPUEa44/d5UZo4u/GD20qTe+6eYm8m0JXkdL
UPhwY55+B+3740kyDnk+uJARBV4k/5jBdBHCMHydY54NT1jgTHk2yLh6qZh9P2wwWG0+AmPDrBHt
uPbSCB4jkT9ETu63euDeXla4NT6FCPrOskJy2OQ8c9yd/4Q8ozFj9L6UG8bW5qrjprXKZ4fCaA+B
yQ42jq3XlQpgsBoxDMDWtwGnRXHG5up9MjxG7s37yJwo4FuUkJPP5WFMpMSXlj7pi6TRrK+tNPYk
B7+J9IxT60APoBqrHMIA57xnNTGN7l6F5vLE8LCcD1W7D0XM+Vuxk4F9HTk+8V/lghRSl7mSDmGm
fueHZIOWcuOGO4wMwjSKiPku455lTDL+6ppUJ8IxL7USuj10RpykZ36HSGEOyK+LEciLJTnyUZyk
MaJu9khIzAysait/TnC7yVCDM9loAvuiqkAWt4/YCUhfatJ917dxdOG1eS81NvjvJIMG4p0FY/DB
yGysiYcCLEyzXzLhg5wPhkMOcfnzFTTvjgYWWmBrM0nVFZN0xdffa0sfiKjoTFvpwAVvn2eFvk07
zqyu6vGygwc62htPkPQrgzMr7RAvE0YxBo8ik0TrvxFoUYPaG0I5XiY6Rzb+CNQxVU4SVF6oxlSL
y2Xig+B0vcl48op+juaXTCoUSGv3y85JBeljZkkxDQqbVf7DbgY+9Gs66TPoPskihwTETIPubyKx
O6HH0ef/1nVJu8RhD5FK10O6A7SWUzBkedoY02Txt7gjwxz9UwOl7LLaFd5hsEnMA55I6PDvyPR8
fpl6w02VU7gaQYQfLfp6nOeOcHGsQ572mbVckaGVVLrU8kvfgQzvDL8lsqxjPx5GdlELD+Gfr04g
4Lcd9hXD32eRL8RkBKV2dfiEi1ZHYTgEeOe8tF1bRWFS2/49Jr9nX78wHEaU8GKvkOUY1qjtpRwf
y2YqLZCVvy5cvwcgulfXVw8X1EsTgQK4srpWbc4ESeRxcAcPq88Xn0IeGllCZT3PIf8fQelqBgjz
0QnqtCxmsYOIh/BF3hib97yUwBNIF4SWETzYPNcmxMLKjUfaFjxn6AJS8GHoFq+97bsQ63xy8jpK
HHEDvmPwgk1dBxioXcmj0hQqbu29kGCANnVwsfzyXcyYtYfniXjXUM1S/Xd4Av48RhTxEpuK7d0f
vd0875+CsBWMs6cgC9oqxCvauVzATxrDJU7/UXEtS2x6gEFEAxGZcyI0W0IVRSZqBlqepY47Ym1l
Jt6HmhN+aV1C2lPXCACyNqPaNigHO+DIodxqAHd0q990G5VIK1fT1uZD98zXLRSGSEJ8fydSDegD
lNhHP+2Ch5Nlsd9VVwEyrfRsT5diinDEPwDX6BVSxlLejXRATlMZM9rcUVD6k3LEFGJ/pzISPrsR
5q2vdxZRejDIZbdFZinwzQ4y2GjwfujzQNALHQkFKCyCo59AwW4I2sjOp/h7ZLCCHkbaxmEC9ejb
YnFNjaweoSOWT0QPRSPpb6uIXsJz2bNcBUcI0BsY9Jx84uHzQlgaiwPZpkf3ikd4wQ8fJx5Ewe2W
qNpre0yAppuSw+Wb2IOy4CkeCHKSvWjYiOSrSVKMvUMy+GMVFQ7ofJsRLYZ6hpMwuoj6uYqkRNT9
Zq2BKxG1wfOPYONV8VUoub0iHjyQRbXvH1cCsrSM69LFW4m4yZaTs0GJ8A+3i26bjTdXn4qySUY4
WRCrBZkmlR6FHnoT867mbuisDA/BUDNdK1xcxO8gxolJxgrF/gcPfxIivh/hYwpDzhMwQbuGJQHM
nKoSkrcIFIQHwHVPGORkHCFUSKmLHuzSqdtFURRmot0U5t/klmXAaf902ACPldhdxJdJfT6Dnqdm
+0Y5i67al7S5zeyx0BGKkDv5j4nGAHoF3bX50CLTME28tGgsRO1SH9HZKOmuXzVJDDTDpZaz8jwJ
GehWBjDrVnRf3ZApnUl3YPdMnbyfTgVdfe9WV7GrO+IyrUnYHdvkr3b7mG5Sdo9K8pw7gbQf5IQX
bFMzdKqMkzmTc9EMTPLI/kp2Q1i8kbouTfGPUZKREVhctSg0TcKs02j+OOslEDYcLaa+XxBJol1a
5czRTNDQFtYv3cZ38lTRxH8iMa1543q8MNODQAzhHQ3H/jVgv09Q4iSkcDAn7wnXZ9ZgOHDN9F5z
aNfhkYplCj51E0vr3TNbBu0+ZP5R+kjO4Z6FkLU6xz0UlJm7jqOAYw1pJDRe8hk/ksW2on1b+wcR
aEzWuSffleF8mD34DkwGJ8VHc3g7cQ8BVg4MeSpK0162msLKzi+O28CUSVgEbFf0PeYdyTXY/Z6l
SZLcARJ++rNAMxZOMFFBZkwCgPbRkxD7H+TWEFlGvRWh+DQKi3/p/UFmc7QKhRP7w5EiifjHdkr/
7j5pQ86CuU/SUOy1eCoqOCjs8csHBierIDt7KzPv/MaK3Y7svS8Fib2cxbAC3G99eyg9H2DwJW+I
l2oXV/3H+tvkTOgQ0I/DIVD0BZJOArfCZDJYHkMMuXfGx15qNhjhk73Tqhb+wqXnMymdbFOWKbtS
IJv4+DbxIODrRhlrU6+950yV1iFnZly3+ApRThVqxlc63SOdILLsJ/pfaWIUqw7XHnAemDoQ2KyT
ZlhFsAU/eCL5cqZzFQOaiTgZ3LNzdoqyXVPyvK9f0Z4VZTV4sH/awqsj1gv+yCmP0HjjYK7vSvsH
CWevAs2zbu4rw0qzg/ne1jYiWWCUjN2uZMfDoruLb6m8wObxImRO6xPppnsD5JJ1AkloReemmq/j
jJnRHHQAchnclDn5p/48XiDUsy/zvGSsG+PmkLxdSC5ozgJg+eFca51O19u0ovbfO6j/L0sJP4Zo
dSPj/DheGvAJimMF8WGpn2VI4z+H8ulaP98xH5fDMXMacmzBBS/Dc0UE6tlpGAtot5sKD4C+l8Fe
3nYJJVwvl/gMTx3iwRzCihpM5f1RZSro8nA6QQg3FuXTECQ/CM9jgBfHeM1s+hvhMJdFn28+fAHr
C/7i/ZcJIiRqcX3gZCl0uMGyPiU4nQxi4m2kJowz22sCLZQnYL4J/GHp3Q0degoaLU4xAFZV2cbC
vhbxaiO0qj5GTQ2aoI8sqt/hhKqi/TgWtUN9g1MHVSgL1Qqv2UFx7LsR7/jNfLiATqim+6HCXf8V
iQUpmtrP3hWOJbkFbk2HV7+2yVhvSa2kl3CvKEyTRNh45Yqb3qLm6eEIlKOl+zHp/K9NzFRYC6Kk
sbZIti4WMRZP04zmu2F4q4B3bmSnsGlQPOrBW2zdlsWxqqEsOl8vCRpIhFBlgJnYDMBTtNpJUr+O
zuhvT08UU2oVbMp16p/vpNl5gQ02ccY58eB7/DnPCOSEHc/MiBS6SGJMGPmkCHTKE2v2xQWxDYyF
hCIhk+xaWhKeFlw7uDaDudHsSJ2VEm3kl4qwoeVfM2DU7Uccdl0U7u/IJzxTSIxaGghPVz6HCngp
BbBNIb0HprJqyqVpNJ67mMjQ+S+zHHsM1nKKy52ax00BV6vwk6ChldpbQCpwZLiVaeDE+bbGrR7+
v1MuEVMeTiC+3aamIwNbJurjFnzWQXBzkJGyWHLbNO4J6+waQgoRDN4etNEEFwJKDB//uUBBd3He
SyT5DaYlaNHVmt92/Wp3lPE6WAdXv7GXeRE2VCJZL3STNtLMkPa8FM5py4AgZqNQ42UGmPLdVSLq
INx3ohb3fzYKJP7K3E+g0nm9qJip27PPmvl3SaW7eXvV1vPRQVnfjQI49gOrvELknwijSP6QIZXZ
A3q3Yk/tXfDWbCEGl+qFymDKoL9kvmFhBMXWqvAn8sOuNi6xigyRLbHo4EIXALKgpObY+2XExetA
1JWbHH3+XuNaS61m0JtTi7W9yPNkbfuIrrJ0FEGP90yCyuOBO55WlYtRCv6fRkQjin+IbTRgO27y
SFkJLR1Su2flaqxW++Od/D2nnRXw+SYyzgelkp8naEXnCKpmD57X6cgD8HTXkwAnlGZPtLgmdJIX
SdKxb9UEwFdeRzf6imYJoFNSijjV/upJiNA57M1uo+P26HJh9/34xpR6wS7p+bECh/5yo8h1EgHs
ooikgdwrg0qTAypE/R1TawY9pQ+uql1nW1G46jMA7AGQ1CShEeS6qOS1ocFrbUnGD9UB8oW++Jxp
kMR6qC/hZKxfJbgou2vMcO8wY20PA+ilo/6fwEkMUvAlkV1adRVNcpR2SoHstLKLTlfE8B5d1eRL
8VCSMLflQC89Zh5Em4vN6PaDDSQN1OLBObFdXagpRIsIsPSMdaukojY0YBzAdLw/EHs3CY2uCoW3
eovG6hMQPSzmi9ELh427WIdt3E1STJzHjRH9klEfjGiR1hEgAO1LbfRiSDQ/k3soAQcz9OrNALxv
v3tQMT1rfxkTjdzB0CyNQ9klHzTO4wNSiVkNihg6u+4QwjbhurmKPV2xpX9icdtkCvqJFRFOvR7f
SEC5qGqI093dRhKjcigcoiCUVATzhVMnkPK8Qb5FHaLpUxSYOSaP3WEV+usf+zZzc4UoOY2mBstB
FqzaZ/GwsRHJQHnAfZMzG5G91mklmlmqyoCAcjsjQx+vHw+AIekxd+jFGbADg+EbWuJ2PqEgsG0Y
YSoWRjvjr6fglRqz9aQNFGU3NZ7Z2aKGAWqu96GzoHn/CAc5umPz1e92CfVHKoOWGfQ8QfzPLV5z
DdPrjxWJ7LINbYG5kGBI+lHd+7vOQxDANs3qhoyd+Up3UedNP0juHYr4QbeQ6HOAhJz21Q7LXDvH
chzjeGYcjsxeI01I6LBqDaH48bhcHr/xonFAzhhk027/5cCCPVfFsOnZlLyxIxcfvbmO9xrqRMCS
qfNmHCQjA0tFoG2RCaZdnRBo4xcQet/BmfGK/vMZOM6GsVMkZawYU9O19TE2AMAiCwdDMk9Yg7vg
QXGpTQLbJDFPnVdN2OHpJZUACfPtZ++pGmVN34PF+PpJtvwwmVp+/oBmP1OJDpuW7C8jTeA1ODZR
PNa0gadczzyL+cTpNZiYIPjet0JEU22ekQGI5MUBBcrTY3gKN5gYbHQBrRPf08cWEeuP/S0TLqS9
O0Oa9Hk5D8g2UBrf/bNHkPI6UVb0w/u1E5gBiGIltS0WTD827Pgz15GYSBGx2G3W+PdkbGO1dEsF
6zK+T4pl77daI9gB9suuN5a4yN+T24HF28hOfeE5YBgzqSq/l2TFOp93RiNEOQN0/LL8lb7iftXv
1Z1r7IBHZ0XsCzReSu4fVUYCEjVTWp2iel25VZOer5262oDQ43KN6OCJbP7DMrBBN6qQ5MK21sG5
5iWuOOKGOhk6+VTjb1JirYnZoIZl33vU5nFMOKTGm+kgrF0kZR+L+/O7r+p8ze6UhjJjlB+KJ4Un
XMMxUCRyP5JPHtxPf4WGWRwb56xVdjhVtGibTW7/cuEVufwn/QEsM84uui0kBlJ+fdfmuPEgV0m+
JpA/x6reKwesloV6XpTscFWN0NM1lW+tRtWQmefmgYGOellP93SkFL4uvSGIDGPdaPTEouGV7hsp
z5CeUeKsIxSrxBMCgGS6n2c+w62QVZwQnlTLJ8UFJroPsHNmqr3xUboYyOdvy3Aeb7nHK3vQ91MX
hNwNtb2BDWBubkbjfVNfY77yx6ed6LzpvpPdMyzelIm0Zb/y6/mMsyHfKSrMwFo5M3cRW3zc71Ba
MygFmJLavzP0EJxu/C+zFbDtVd8vn/Yv2sJa50t4lQfDSsXabN3R4Fjf3c6PavdSdUHBCbS5GIT/
3eD+bE15nzGitzsyDxsiX8F/ZMPDk1FrMIb24bZ3TMFV9jgoLggbH+7cZW1hbLZE4oY/Q7D8GBMb
01cl4hSFoQVlfmQfbW90RlqjtwpAjN9uPkkVBElYxaNM057xxf/qbHvXjVV+EnicHI1qdBPOl7ES
1cnxW3+knm8lpDPA+CutmTrCNWfAbqRJHRRXsLmAV4AamcDUaxoXtA02bCQ3dWIsYx+mtT11cy2P
GIBybN2HrCOSpmElSchvud7sVOyqTFUlMsKK2X914H8RAfGMM4BRu7hvWk/yOYOveULfV+mniByk
19GLke+6E31P8lFH/zDSJaeSTsLJRYsIe/jZa40HKoCxu0qQ3Iq7JP2HPg6sZD60w0snMxB4IAf9
fSlHZbYcfyywRDxqxMWm5+JZat/uaT/Zgr4L+uVIK9iAsGupJoy+kA0tZWSZrz3k5DpJVzJIO1l0
nXDiNcRoIf0Do1/VYlUdmIjXJB1tRvpF4NJWyTjeahgrRHmReTqV23t5PWK6YJhB02rI0oL1D1Ml
1pQStGFz+CtG8X9iYdrVXapsRCdrswfIB4RBfkmnH7HTiZNToijWT7z5w9QiT5aLsvDZdtFTz95n
6IiX5K1JHwVbiRDI9zRoX1GVjrtO7cdR723zTHdPGZI3aPoEwMdN2lVB47trnv9D6vyhnk6kqVLf
wk5lS71YD2WpVl8ec6gPaGZBOjZi6j4aEZDXgwbnzI6Cox9qP5yAEgP7tfEh/Rp1zWm5ueG3yk2m
zGAOm4X+yaLO2T9bRKaouYNhSBIWJxDO7ytsCgxxDHbhFU8LE+QPKZZUujBg9blOkCMlAyd2uwU6
wIgQQdQhTNO1bkjCiO/uekec++ELgklxm5S8p2uOSlGR/oNSyMHMfRTvqZWTdQjRdpp4HYGozdc7
m+kxxNaRgPSd7JUoy1GZb8yqDZAZScbB/q7uqiBLZyahInjHNkkMO7ZRB4F8mhkahxH8HOz3AkSr
m7TaaSgrbgUd87pVe/utIPUd2oWKljBQaSW95oT/RnG1DLO/pBIkh9pc9hrvaIeSzOXnYVk8UG2w
tG+ipnkrszLnku3I6HysjROB/bZbDan0DvgRZ8o11SbH+tUWusvFaACqUpvVJo7MMI4R5UM9eMvV
UX9IyViQPoyiUzkihHpTTEbdzJy5OP9DiTKmbJvshS3LKQbYEu7H6m0EKHSI8iN89DpMSnpG+vmI
28md4IiWD2AyFOLu+9F7MoHOvtE9Ye/54KSpLZh2Tmj5bokLEbhCUKOgEhaQpm8BnXey6w85Tpkj
1La1xEuPHTsj+nB3ByC/CRH2cNH8Xyj+GpRF/nlk74SgdMt4pBBGnxY8eYE0NIsWlA5tlpGcEUIf
5ieBjQscnGLr5vY+DE0xwbqxa1ebIptd1xLj+DTbkjoo8OUCve+keWV+0EWrw19mVloYf/yyTJJQ
HYxhoZbITrNVuGjdis+fd2jKGYyVT3ZdeVHNj+EJOEdPelqf4vkVfC9nUCCqCqJQ+RLHee0gmFyr
QGmt1f2DH0t+Xep7N490EYmRenjPlM8H+nRLcLRC1yuKqBipobdmgGOR1fhSWPjVxur/M9b02RGL
feSzmS81ad6p4EiSxFssLeP9Q9q3yQ3EBqo356fL8MBUQAEnHBkZNPFvHq/JEz6N9sTbtwKeiRSp
mmwod1V2pnFbFHvELDFCO8uJlpa+/fjoWQsN17HKpf0+uWsOFh/1L6QlnTlO2ocygGARRXxXD7wK
2i4RYLZ43Th/j0R1Xu39pUdD1ge/XrkVN3pIrqIworBOn9NHNlXFEmhoMuOpzA467iVcHj9T4Q2d
ii94t0wzPUzpJ5oFoQxVt2BjOijRsnVfK0cQ/yi7zb9HKt4t8RUMwtXOQCzO6Zi8tMVQsjwQqPxo
qxpNEuVH0git2q9iXbhD9h0wtljU299BxDApIwVZNu29vqduzkYOCQbT0quZtKNmaBKd2y58BX7S
4GJbu2Xa/1cLOdiqym7rHHZ2kizQ/BeJEQtjcWvS2gkIYYBocfxjA/nMdbh/E0GETgXeAnxMWnO8
DBgxGgEr/TnM5E6A6b5Yes9ivIJ2q0/ji+hHgNYRWZSyXMHXk941cGYI+y0cY7Cp09XxA4eg4KBU
2C4DZjB1AyGaN9r+cv5hGe83j3k/VTbAESOXJ5RFegwOLqog2aUs+vJ0xWaFzUyF+4OM0DMc6cZ6
/re+Vjz0+9SocxoQKHdSME6r5kqyhywjaQEacp3NNVQSj0TCy+S6y1JZ3Nz9DkyzOh7g5c2WUwJV
f2t4eoR/8SoVu0HnlwzB6O1eZ8YSdF87b13OER7aIEi2ITAKfNgGImKRLR1fDGnJUZRudlHaadkm
rpxueCmaS0jUgFUQqgPkCUHSOh94YF+9YIMC3F58TQc8N4t+pHAAzcA5Q2w5Q+OzMc/ShTjc8MQM
xDpUEr0zR99d1VrhQa42Sm6+f8aklxHUc106WKVIC49d1R9tBdwp3oOyG5F2SVXVDpjh2/k/HdEJ
B5+rsShRMnXmlx1c3suK/K23VrYH3adOWtI83a3yCl3MPqWlt5KlN6fcpgtolFedtmXN9VJ701ci
ss+c4a9APZem8AJhRPUwBIXszaNwGdX8LGfJk1CdA8PA3A33VAmQGdninNq+XRxBX0PfdCmZSYKX
/Qsiq2HLiSCLnxKcVNleQudIoPrbjLPoh8CdXimt8rOgYXR+aWsSU8vDcun6DQ8XmejBnKagRdey
fsR8+O7ZZTSxEZe2j0KThK9Zqb9+GpKuE+Fk6w/XbiwKns1r4NnztK29Px/5xARcmxTEq1b8s4nE
sYt5Wbx+rBTT0wDRFPjaC5lKylzGyc6olUwBLDhJNEoL5G8wfo23jMF3u7eNiuktp6PABmLqQZrY
MBo0rOgpC/5KmbQslCs0IkDl/EORoFbt9mx9PVaIPI6g7/ONhSeMWdHLbhvqnQbaZeFawRDzJkHC
ssopB1qNNULPuhHUsauBUOkIysCdPErwNlj0AQNtStijQKrqMCh5Ob3EKDTr4+u2U4kyrmDtbeFx
xcKg/ffEWb0wfGv5nHYoEZBJoQP+MT/gYjsG/7KlKLha3c8hZI4yEi+BZL7+/VWBgPVAHoFWlb13
cVj++1GhCA5r2n2vrV+OCE4bA+IhMU9dYk4OH2rFB0BXSnqXgtZ9W8T3Ng+mUrYmx05saVn6CPZF
rsnzUJYhtD4isVCh0OKKRKzgnM/+YwyWGuGPIrbE3sYMBLAvz7fepcN63+BLK/LOeizeJKb0JwKh
zXHoIxi4U3rbyCLXjArtYcBWZ5E4bibq7tp6Ft8/0QxiEeLTvo0Hf7hZKPxud3MhFOuTDZAz0IUx
YgrdDmdJtg8eUdWXEWA5kRSJxQabPiorQKKWPn9wBLdbsw1Is4hO6XjoYjjuPgaQBFKhyfuXFArn
E4LOtiLzrLV7WDxaYmVdQqs8nNhgBjWOuOBH2lNnExIOPNjv85ZqiQ6HJd+fw6AUO33UQA4EnMqV
wOkTac116HhdtUN3+Slbykkz1/Tuu9jC+bjY2Y19tAdS9tBlMhT5vpw9OcnqMIngiEvArS0TOhCO
ASRjTsaRPMAPUSw2mM+DgT/vbhNmeCGC/671tp/s3M0wI8X7MSBHwk6W6cuni5MFQxVyI95lXJmY
3AHiRduKqdNFZLlf883M0plTQ0TPJaz1zcR7sDxc2efHkNPPlRnco96uUEkHW5dv8Hnb4CVjk8Xl
OvkLNFXgVewVX7IX0uNw1moGkBs36LVQXTum7GneHuzLqiWSiyejKqzLRhe2eUUgjAL9IMpqBUFq
ZzzZDC/9T+3eUYzGrNxegEUG5440byo5jIqihnQKtkk9VBLlPun7+aYT02H6C+y7MNsg0MUUS+6h
Kq2rNkIFVXogCuEI900QrV7TA3QaPeqcXD+8eyAssOUxCwr5+Z4/k3T24BADolpK1T7G4LSnQAnM
iJmk80IeYcGIDerWWsc/9grTFkezo+BwhnF5e8ViT941X1RArC7eSl1uvKOv097nCTvGe8oS4xQW
sA3qNB+t8gqX2rZvXVqsk9TZRN4L768SWBVcxKVmAKBn7EWM+2jMNg4QLPwDlpbdtu0qBzQc18hv
MRfqZhc17PhEL9mC9NHOUnfSRshlBwVWLrxMByVVSh2Gkq9G0cFQMolWeNjDVPxnY9wiYyn3MDf2
asLlFNEntvg5YnUteBO+asCgFliPzn3FcmIPhwT9VZfxIOUQWezoehLYfHBSjF0VXPJZwP+gHDAs
nPsn9d5RPUsctE6Or9N7g6XF/B9oYe6r2TALoGhJ+icdm13zY77ZRNeEa5L4drdvsEFqd1CMNY7C
54AX8rkDmLNSJxdvR/ZnWqio4m0qgft6XNv/csYhFpCCW6ghnpOqRWSHCADwDkgNW0zhbpY8zGjX
P9oghcupjid1qgSnm+rJU2uxZkzLn1CVhmHhU4PZs82deovhRxI565QcZsleWYv1VlnjmMcoojCI
vTNf7U6TO+2PbCmfGJ5aPQKFSo2J1zc6kpydWNZnUW9imyS5cGs1NgL4BINkj34fPV0GvIgYA0X5
pa1UwiJaKQNJzO3f8iN431I8nz25JIdQb8f5jYIKeNNz4h1Zi9blw3Zy2pok8VrehSON8IJa6Apq
RPukiu0og+Wd4jAfjyyTYQlsC4GakMfwIFX1/TNmv6mi5ogyRZefe9SZdX3c08tygPCa8AXiDWH6
wwgGxV48rvSNK7wGhIBPPewsnmJaXDbvbSR7k3oeRgxu48NlOyibleYVaduJToTR8jpCchvpnzkw
AW1p3IZnOJ0r77074lMuig8nC4Q+vsY0ybFgjaIvDMLA1O89Y/lAc7HLHrzktE38+iHfDH9D4+vE
huHO2sEvZoW+qliVRLp0mg22k9tN+k3PAGmSX4POVWTsTTq05opokXY97Apj4O3xKe+j+ggBYQ72
laEE73neuSRO74jk4bUbJ0gaAQ8qDoNFVfwvTWx920mDPnradv7eW7z2fGCVHULnPF9pY5aIE3oH
xYV9MGUZH8qlPS1Fb5Gq8bUpD9rXb5NpV1wd6smeCc4Oe5L+5FKCxWLfWsBGhKh8RQGhsMSvFxtQ
4nSV00pFUXTZimWtopapR2RASC/SBhaTcgU14c4E0sKjrRNOK2rQ3z/P/8JsMDj33QUyZtGJy5Vy
Dly8Ltheovc/q5zz/1e6CUhsaSiGoVwimqpiCjKgGcRzBptVHQk7GH7jwPB6KHAdvtG/9I6OWdXB
sZdSnbRtevpyMCyELV8GUV6QPfPDwIceG33Ss93XIJjS9NBBBvQVsSczKp9dJkQOXgfv+LllTZBJ
XSLI+H4BVA3v3bY/M7bK0O7cprYI5THViGyRh4WaMGk3UVvyzZ308QlTk483tuLs69C0QT9M9E3Z
14wLsrqvwhKSSRD+71yjhv8We4jp5emawa3dYXlh1bvuTe1V+eaIiVFXRVEEQ9tT3vJ/cAH97P2K
Ys05qlH/SvSQzjBj9tJr0S/5WU1/e2+wVu9yNSkvOqo+/t4bMm6PXpse1HrVTF74HgqeSxNqHcp8
pjLh7FdSCxriE5hKXA7EL5PDMnp99wXPOs0GHnQvtjjrCSD7lMCERBUBNvbG0c58QuhweBZplTHI
vvWN817cpr2xjR85nY3E5UIaQ+SVGu3LlSvtrKQCXyLiTHySOJBGiGtcnAbu9nmpnPEemUgzVryM
MO+5KOyHQwNcPoPBB8+jGioFyozZJNTJwOrbQQYvXf/ZYr44PKsr+4v3ai3zUB1EpC2O09SH112O
f3rRkSkGYkWNpTYZbn39iChJK+db4GtZrZ6Nx67JIkl/0BeJv1l/wfklNG6dKVs2vwjfga92IZ/Z
j2+m8o1heaG3PDpoUFi97oZ7uvkXMtQdd89PrB3jc0OLe+ic/CZxh+LmXPQQHXCQGCTN5wIyGFaD
Nj2HCEOFG3krUzff3kxiAkzO4yFt0SJn9G9VfCpfoHuSdb5+krwrdRs18gvnd7aganDHEYHGYn4O
rJlJxtJ8CACxNAVC/EHT3TaS9LW3APg3pgGfYq31hibhWACyS00J2Va7x9TsmSGww60DmHgEU5Sf
XM2uuqUkLMC7hpf3CwqmHt8+EtqqAQX90IAG4sjrz7baAF3Dx54nHhyJUdQFzTkaVAeCu4/Mv2ix
MsnrXkRxkorMCys8Jxq6xCkXWf/w/gd14mHXrbVUmmQUuVpxwgws/XkpHAs7h0KcnZmF3VrJ6pZz
dGNWm9IpzDjTbLjmlOb5VUGFE/6fBw5nW+9LyIsLj3/MyEMSb7Zoq7eZ45Rm9Umcp97cFlh19ilw
XFfFj1r+4p8a/Oo0Ycl7V+4ZpIkVFLqNipbEwtkcMEa5Ce8DmicmOEq/1hvK3Hd9ez/54cDPwFdb
clWrzZ+ceu53iDeScFhrRGTZ9YtuUBQg+yPyGmhtwViUPTpoyD+ySQG5AXGhBLA7EjfoP27beuTQ
D2Fi9x/JFwBh4NJ+mrPx5OEjHWbSC/mUmdUlrtvpgG/+saC96KRwYFNBUbwvEuGKUuNcyyeeurXW
nmf5seS0xcg0mP3i9odAejkgNPOaqeG7BiIY8ID59QzLH9R5MrSDK1E9hfl/KeO0oHsgsD5no62c
yTSlkpYJDtMH8psb5dcvJzxE+nkUmnzm6klXtBqaWwzdNwueijsPXd07SU74v7qat/INidn0V0O6
yMiDcYZOlAgwf7QB+HsKV4GqEHC8l9WhsnJT9euYgtkSlBUW7Q7B6tFZCPcqNVGPqzmG01cWk7/9
CnwygLEm9PzHISbfiEN9f0hpV5tEcB2QkT94EZgEr34dlHriRgXQ5PvHwUqRQ5OfQ9JTofIDdM8o
XmTZuAe5UEdReoD/+6ksyIvHu/iK3elyNE56qq73l21WaTqczPmnLjfCDmlPxdShPabVzK/XiTjJ
ztjtW2PBTLR2TJPp/+PS1gLFhX0zrv4a1TNMF+BrCIRVmbbFMQECNX9aPAcovjBtOeKsQoxLIhtW
UgvYDzaNOqnIszC+g4TrBJA2fsoxlbV1FpBuQM2j73aRWNDwRZQ2ULevbcJ1OXQM/cjhQ6GYB/OB
DXbipENS5j4043nDGWLKgQG1iPQEG6m2LADEEOB6BAypZ5rsv7IXI9jfZe8OUp90jHoriaZhPur9
kIiN7d9Z6bmfiMYKr7bBGO1A3zWZSxA3C3U68EiqnJQ+vzOyE6MgjqNCsS8YGPKaiAkZddFQKxOD
r330KKaoeDnKeT4Gpfb75XzGnAikOqTkSAxgbBGGdsIFzSI4EDbuSQxM5RhPl0XZy48mwVcyENr4
JDB61BuQn9NbFO2IC2BPmz76nwK+HZ5yK+JU/4JL/B5zpBiE0c/CE5zeXwJoWygu7+Wu3AwC3Z/x
cySuJ9izJPqhwWLBqEoKj6LtxlcYFyUuSlNlEMYiUqaKcqBcnjO+lKITfxE619PuTJOyXOj1/qRA
QcPxma89HF6B3/xuFLWbVNBO84a247RplOTKq6fP3FHzH34qcKnE4LpiKCKY+v7YO0FW98FQmIX9
hUzMfUjvuwnss8Tn7CI6i9+u6moVJjCxR/IBO9wcllvZu0ljTwrxqx7aSjWOoQJ9ZB/4nbZDPdCU
NhWA0fU0i83KbH/c8g/bRixzmGCvZE+92UJWApVBpnUNUu7kMW+wqRasLuzP7DJtMba4p5+JgKe7
G5BS3T7dsJrBfpjles/gzSFoziLnS+EHN2GYTl+svlW5aN/4FsuCpK3dFXuvLHvP7Nebiz5nZmSz
wmgb4UwA1crom4uC1TUwSiz2VMsl36FEtzHVGlls1gqbRBBdZJSkziQYKUFDE+cC75yjsWvvuFua
nlViUFRmSJYjI5cZYMNV2O5t7LMLz1AopgNdjt1oxMoWba8l0WTbZoGoYFL5sCvA68Q4Uv/NdnS1
et/d608oLchf3UW/rWILSUNbR74/B3GbDLKIUbLPrAv+wRhfXSdyu1sVdJ5Stsz+TY0XxLOIy3Lz
86U/k+dF0W4CojMXvtGNcfIuWy9OccpOdAzY+4U9kgY7yDjJksr1/tep2FOp4I7lFJr7khNDjSvO
9WNNV+UJoGIwqMZJlZbvHGmzax+UPU4vK9+jb+KFeT+sx4dRKOS39Acm7WFeSiBP59bvsyOW7V9z
Rih95i2B1jIDX0d+Gjma90hLc/eYe/k5itTBiucFuic1EYcgBS3bgkhNKOyclH3iyKB6xxTdgP2n
vz0asB8CrP0XfJA/fzJaxo6/V7cXGdcGvezL7LLK9Zr7v1caPP8gwpqNLkSkSey56jDQ5jeggiiw
tPgKXuCbZKL1TGPWY3wrXJowDPzq7Uoixw/eV9+JUZl+6sPj31Xo/AZu6CV8QgoVwmoZ67ZfzkNZ
HzrjffHjmSndi9hvD/MCwy1H9oiJqB1AQizX0mgKIO6TQ/h/4pSoBizBeF3dVq2qJi8ZfgUeP6+N
zAHOV/kQoK4m3ngfkRkVVNERS34potueFvwcQP1SOVaMvymSacOqO7t34Fl4l6b7TkV4isrI/Kzf
aOTRQA6QTHiVP7JgMyozIVZLCf6Bjcs7sRLNhatwUqym4tFJ+q8KRl3yfnKe1ZRetTsMwGCH/w4V
AahvTEjQT4DtzE8itt06vvp5EIHJsmM6kcIybLtAoprREWLbjukPPpaVyYOz3kBHHfJCBGdgxll8
DLEwHDWw1R3CkPnmX2fWQo79M7ivI6oTG7aoIDXvDtK2ibaSgTHxUHzXlOw7A97qAkqh3nhQ3Ob5
jeI+mraCGoF1Ex7kcle9kOtWKmBaBnQoPm86YaSUeY9TFgTlnSUdqS7tL1zlDtPr7YvBbDHnAUCn
GcFJdpIXu7Y3mHj3JuLgSP9fUgkxJtNjcF/3hF7W6P1lNWZumgbD3PlN1vgB5jSmMjrjBiYOR55a
9RdyauBTgn9FX0JtlRhM/ROpHObL+wh2i5wGcfQ/9YG3pEvrj9Iec3WzCJ9Nkk35uXLAtgHVzOiB
JdAN+rLTSJJwF695Zb478+dm9Te++4+KlGEXTIvJYYcMOMi0ULSyFebkkruqQqKjaRQnp6AWcWco
5VKDOP3m+4s3Kojc0K/k/1xM+cOds5yR8B0/kkrI9Ee2Q8NLuluSSl8lJiL6HnBBr2EXOWE55sG9
TQylrkZXaXDVuYq3ygwUvX97pVLMVBJVcfjJydDBYBotTMLjTiEebvgcUrD5haeCWfngjrlsK7vk
L9MNEb/q0AW6rpOuMeF+e2p4/yL7AAA2PX5UoAhvx3K5+4XyX2FH+BjpS8G8GwrEYkTNBuhZW83X
mE5kDcMFyjRfvM6cVeYNuLbqpc+CamBPmnrTF4UxWDfgXIYHsNWBGp0EAB01hv3kpQMGoAuJp3hI
kBzqZqeJGInAK6ksYuX4BvHZvXBJCT9BpMJJ44JdiCzhcL5XFjTqsOtMRAwsKe4vYgWYesgr/UuN
xXEKj6WR7sOvcT6DtxApicv3fzv7wx9JnN4hMBcybni60Msrl6u01ea4JsroeKRun4VgdR8mkmQs
EdPQAADrNTzHD4S1J7tT3DEw4aqle2FLJuQxKmQkymr47hQAeoJa4XtIuBq5EqI7V/Jv9GTJLEDP
3lnzmEDex/M3I7FcrdUNpXwgis80HDfWKQ+SeN51evBP1A7i0DXI43Lm5ftF4p3VrUJKs016S3zN
woIwk7/hyfWD1biv+Im+40YMf1JSJ8PUSvtHvRJngWdzY0G+ZpPd2Y0vEjey1kH7vCO6Mp98Jff9
JZ4ZCRQf3S1G+scEhjwycr4JO4BozYQdtiuCFlIykBCxPRUDjv7tKou96eTaStSpUdBn/CncrjeE
QSHfyAwHZ8lWXKKfzHDSmAbt46zxDcQc0ZlJE1ooBwOv8Cg6P0UvOVMc8XCqjd2c/li19b0kXPY+
+7zT9RbTkXjXhMaoxOycksq19UkfGYfzDSofs3f/D56liyeP9eSwqhvYOm5396oVZJR2UgOSaeN7
tjhwbQBLULXjQIfxZ+JjXKA74M5/iN3MZFfaCPw9f4/0zexKQk430PGLJpsQ2dNyS7Pss4/ssU06
/l1buwveruOSkmB4RIi3g/0jC4zH6oE741X8+omrXs4j44dbb5KJrmH5jXwQZW/yMecvSzMYxj4i
ZiGP2nCMAq3YVhcBXrePcJqRqYIF6j6EJ1j/VE5JmZhz8wq/F0IRXlzs4Boh+im0TdZVpZLY1bWZ
UpsOMWLts6Eu5gIOL/FWbYu0OsFBrnUB2I7lxXnS94ZveoiQQ9c09Hpfp0CBrty0D678uYIExEdm
zlAFz2gM70zHjz07MFaFRUHKIS1XrA/BP2Wv8m9W+IYVCxG/wBVm2RAD8Y8APWWmt8a44bMSaLBa
eoLNBtDK5NSP4Qz9143HsZFOMZ0XN8Nkeb6qHLf5hZ5fN5IcwiphSgxkq7XHNpXtccVtLQYBEO8x
QtQWw9zDeSMlJFAC3ToEAh3atmFoH8Gec/g1YzlMukSPIHB7NibYCu5kSlyDuyJ+yK5wb31PSolT
HgFyvLfy0+ZhmKPwjoQ6ru9/DlPHUTaNrnvKeLs210/WUxuh7TawuASllOEWxbmyUe5kidFk8URh
mh/5qjfZqwG3ZWJ7D3z8tQBctTHz5zlAvqsIw9gXFSOBTQi0UeKDy1VctvxNREmyJ/gGQG6FjVr5
we/DwBQ/oV38tC+2Q7Ub5kFxKjCGMSNVp45wK1ndZOtX9YKPnRjpu3I7cxcvepq3fRbzkgA+GK5D
ry3JC3MxJoEyZw03K6rniv+mvC27vEXu7TemliOChe03LoqYXrU8Mb171x75Hguhlg/XfiC4L8XG
k5bcRgQ4JNhSHulBqpaqCfTBFQdRr+hx+RqUpdJJLWGI/r+Nwe4CI/AFPaZxGP/DGPKiv9DeGTyf
NS1HRCXnevjJvyMlm3Et/eiA+CjEFQV7xdji/l0uYOdW7AW52PBk2if6XYBSXVSkaJ51elpcENAv
7Ts0BbFL1TGX72676RIKHV7nbBG4YTQNMlsQ87TzAGqb29ZaolDdsGSjl8XuVhnuBgvNN2IfXiZc
VhMatkdJneeZ6yfkz+Foh/ftecJeJKVGs3m2MPHNdmL1YA5TQLRkGcR3cla6GlfLm5LahN8iIUib
kJK+YrD3zzi2zWBEilTIBUcYpDR/o6vWEzFlEJle/Ea5C0ajye/uaqKGG6DUFsxn9Zd40bJKwS8k
3lo9tgFRObG4LggLhOKlmjCXuFU5J4S3F7LIr6e2WDgE/DxqnWwl9Pl9tq5tW89Pt5yGfboYhoS0
f5Vh6mssDyBm9eIKtuBmA7T+C5CeVvbAkMhaoIfFFShQs8mJxhOMHLU5+E0AuYmStRXibK0xfkoD
4f08P8qdgjj0ndgfYDjqL+klv7toiOAX66oKyGDx00wTPAiIv1l/o6MyTECYq0RqelqqzKyMYlH6
d5KjoyUGprWeSSJwq21A4nh41MgqNpuuevbMFJxqR5iE9NlP/xeLJWV3+6WvD3AcuVr1zaOK/xjY
VOztiPnUFvvn9Qod5asOqe9u/mC2B8ETZCk0eSn+fc7Tona2h28W1cnCx+M/WbVJ6I+hwRgw50dQ
ECsfMULJrp01Pm35IT0U41LLbziIe6t6L2nUeXZAgR5SDlu+BXb94QGX6qfdKuEibViDAosP+iLE
QPFqxXcptJW1Mn3KKu4j3SGzLOKHOzfB6j5mWqsl+XbRG9WIvgn/rVVrJin9IQ5TDcJf78vL3S1U
VTlijvkSMGQEuaoRyAa9TJhkkWFszaEq9eh7Zw0EPBy3+ZmFkhQVRdBsEemXyyTh2lfxJpYxDNSZ
mSwxiywQSUCRZYC52pbuyi4X5uBwNfteE7WCrJdVGrjZuUMOYe7yY6LPWrgBhIlzwOVr38zOTR3e
fQQO6yIAJJvoXRp73fJLm8owCYEifwyNOJa+S87T35rjyjnwCtOM6Z71PuLRcV1niV9fw7ed72rt
oUJUhjCgrJBP+mJwEU/FaODk1Hhb03fCEXQ7dgqh/XA2PGWciOcSUwCwBQEihRa7PzJIOPo199Zf
EQZLCf1dHWLUlqJObxyFoZKtApGDRSulI0WwIuu1MJUX5DE/Fy3utRn7jHdztkN9GTn5g3jxneEm
vmDrm+/3iHktIeHh2yNx4LW/ev8pkFGiDvb/sdjcPGWp/ArbGg2GKYeARbtjVabvpemnHFW3R7mt
5mnZHG/2F4rgA8lOdkrj9eoaNvtaxqg2Tn+bNlO2m/sv6Y0qjaUbSW/yAWh97D/arbFf8BDYmsLh
FYCM3mBM0BffwEL9Ca9VCjj3iuIGanQL+Bd6hrc1P3IlTgLsAOYidUlfPg09eOnQJOW83vmcBQbz
UeGnmEzRbzfXbGPZYD0iiKahNRdmUZu4K6ukuusJqXTPQREjh6vfuB5lnJO9aUd9ItV9yllxknKE
3qmS9zPPKYmU2BltpQ0SoO5hA6v6K+BmjlROWQ0OOSZ/Q4DHp+q6fpaxM+oYX0Zp4HNg2f1TDyuo
Os8ia0sv0jtSCX4ZDQEPa9wp0cZg/CYE76YYKYXBEUR6dszg846ehraJX1PCAcdUPAuBjZtRcy8H
FFO/ZZu4gMbvYpyn5zYP8NbOooNFq3A0oir/L5Duc0tendCF2fk/SiUJYySNWCAVc4cIFH8RAN+N
hPXFpGI+2s8fVFMH06357GfWyTyYCe0JpZBWPltkWkqGRHpu3bdB+3uegYOMFrRAC2DssNKlptzz
Q1MmvbNAbKn7rWhvwK5SBjQrHOQ9t/b9e4VSXiBpSfQxmHbqF8LRa/hbWaohnng37KCmxuQmgV2I
Jsv7mV6GvDpaG+ZV/pYLT0qRYoCzvUCkNNciKCEA1pAHRrfCLyyH4sX/iYPMgF1XC8gJSvC3vznJ
/FzyQMVl+H+qRVEGIc5poCiRVYlpxAsOOBbLMFpYFgjfTkTx+lLTF6OaRx2rpL9V+L2nvi/pPNdN
7UJKwmv5i0Mj8V6dmEdw1bcsFLSRW1YCm5sqiKcDIwZstpGnteeivQojvkSBTmNHFHM+4boRqU2G
fdW7saCjijeLagkEFhUshfufGMudEXLxmLG3UZijvh023qztssB9rDJYWEwKBjDu8ThVmZ2HTT++
begv9XwLN5Z3mYWaVWy3wnuFW8IK9E2VB928zDqXM7GhWzXi7liVj+De8SPyxAphB9OEsGlIwtbt
sbDGcKm6DR/0SzSc1pR8i3xTzz4XmxE89MVs4DULUJ9Kp/H06zR1sgJzOjyaR2c1ziAxvBzvCViI
FROqoTBVYR10Mq/6i01PlqPhRcNMh0EojWgW9bafk7BZbBeXJMIgN99tDAj0pRuFwSnUwfHPDJgv
Dh3Fpstg4W+3b0uQ/RcLLr68xY4OTQVio8BLVDF5DsivvrDF8WKaXOoXT5lWV2WVAicefYaXuRIu
mSYJ9+2rVIBuCyc7Wl7Z4B8/AuZ8pEsjlYrtVs5OO6RUfYxazWVOE9HokRWEaqH4lg2VeNRa5QOA
ussD4zD49DR5Isojk13gFgpL4N9NiTf7QC7XyS9HfbUwLdigRpD6cF2WXP/7E76rmlYnkd2JioxU
lrIz7h3gwE+7euSsPTpU+szOiANTKdEGR+nfayM0I8+CFdeSf9LnYOvXLQfxv6Nqn5qBSOMDilha
BOuJdXv9hFQQl8DVOvnhFYt/QmdUY7y3YvRcFH2Zlobd3A98PRiaJ+SDHe+ifnSSV5m0x5E9UpEU
rYf7F3+X1RYLAfaaEgdsL8meQ4yP6JPYdbJXb7JXv+1DW5xpUp1KmSFpywO8IGqG4aMCZapiaQNj
Up9bAaO73yFTU9cRueTPWzGm9XGrVPWOGv4ndDlh2csIsF9djJREHgUVk2Df+k10Y4SmOtkonDgq
DW2Fy7dHPsi6ehQQRZCngmiuXJ18LnpyZyZDB5OCqZBRtDb3Zzth92df3QeMB2QqZHr6+YE14SED
FTxPeq28uURH4h73vTd4ZuzoSGqXdFKprU+QeV5edBdglWNMs9WKadZ+CwcIpChdn++so89eKoqP
YWz7aJ/ebxN6f0dMeXuxd0IbSEikV6PkWydBA2/ipO7ccN86/zM0ZFffJKOls+94KKDIEObmrtSV
4MPTMsYw5HLRUhdNVI7a51eWfOxCYFIgUKD6yn4R7kugXVwin5IDnTcRIxXCTWTOovFuGuK8Clzl
f546ZEYEmhlq4iuMu8kBtcMpx7A/HWt2wKAAoyVZ6de/2+UB5I1mQoIe9iEuyUH5Ka/FxQqUeBfN
ZHTGTxiDtKXbGPgdmBveBdvMLuvN5njzR4h3PeGy1WKjBuPOsqeQ8qFUpyMys/vYYyZQ9Gh3PHBz
k2AQO1pk6DdHpPaZGlqmMQ55qOU3R2WusUH7xfatITzj9yXdeFU1eoP6ztQcFTasURAKJjxmd8eU
dDQf4f1tvuPqkBMdzGqZOp3QIF+JwCpGxoPvr9KPQ9h50JpHrUUGfpuU79//lLzUmrf08Qt5gdrI
dJoyK6Na/bMrs01J9bOsnupX5ceFAHyaPlJ5icn+7Bn3BpS/RE5xp1031GaryVXd+m/oGhxPA8ut
FMb/v7aURcM5GIvtky3sK5Ctr4kQJqijQi2nn6heoDS1aEm9nq4anOF9iotWCSPcDN077fs9P5ZU
6bPBq0QqcfZFNUXQBh2BMPuVJc7TL/oc5yXZFgSRmSKaZkAz5gmU9v6UBqRQNCDvSx+pdkRAYa4X
nm4Fb7fES4okBsqoFscKTocHzsHQm5O+buRH5STJA75XggcOrdNEw/mBM9y/JK/BSqx4ploDBSml
cqAu3pxWP2EwytEjkrAjxPL17RT5X6vc2g0+Z6krtLWUowkudtUiNnBU/V0DZdf87ZOTrC178IR0
X6tGCn5ujwujr8LYQ1JwU+SQkvTBvwTpOJ4IMQ5nygC7cYzpn2g/pCDBcx0+3Ov860rSihkXpuh0
DuRD0IfSJSPhowcDaepP0UT+qML99vJHeSD+Dnk9leo80Pc9gajlzXQlSuKKdwgNleS20788NkDr
cSnikZwMt1PsQqzNKiATgxfH8VjM2Z38IfjPuaAOWwN18oECWP8SzLalN0wyN1R7XCgTrT+S/JR+
fX8knNO5Xfu8mUhQOa2wHkYg/se5pmwXw6zs5rr/jMc3vrv7+MlCfUcbIoCFR/cCSuPuopxB/GWs
HS2ngBPnLoidsPikWA8MdX2b1TvnZaS+rRPBBw2qv3JtUgw2N/ncWeeo/b/qc+qy1LWob8zZ2k4d
j+Hsxgn9ae9oVmjAbuhjhNJWMiwK5aSRI3+D5doRgf3bFH0ZtEjR7mHR1jJuE69VpI+Q05O1k3Jb
LuuCCk8uzzbVNRZwhb0YRNjWNeGsbVCUk2FczmHbuj0PuvsYHoHcwL84GVaKkk0U7bE1TrPNn/cl
7CzBu8bDvkf7iSVKnLa5Hf3Vp17NOT0tyqH+ANhSWaGGsPSPbUNDKKegjLrtq0jClsOLndcxcFs/
QNMWGOiyl/BfY8CzRVGmAb4SQBx3P6aR+E1xuqIKi30pq1XIKMSf+lUi5Uw6HEZwkbQhRPgn+ByW
z7/qr6EYYdT1Zgcpcz9Qk44EItqaKzIK7FOqFWhf0bRKS20y8Yh0aCgyvSuQAZpfiZyaKCuxpcyA
b/cRDPWZJf1p+ZZoQY3fmIjYX35uHoFut3O3fElasomDN2ODQfeyITZq2TlazOoTCkBKQ7gdrZjz
EXZM0PYYVbmzLYhLSP/2OUNLCrbMQIIBHPjzGnFHwtKP2qtjzdY2v+E++VLrpTTeA4NMPzoBXSbQ
/sLCdcHmOXt189kbUtYm5DAZ5hynyB2hfB4/IS56L7m9fPnb/497hdOtEVfpOL3MollhrHxQYToo
qGBJbK1EM9iyErzjBvc40kxet6eeH8zwrn8HvWWBOrgCxGvIvZhErY10DI5KVBPteQuGGMqpx7Wy
B/8jfvnFjHk+c497WnB3pY664dBypUDt9bp0SUDdVv/jVsX+iOZihmCCbKd5SuguQwJwttSDTDFV
TBn26l1o5S8soy+S3urIOBrLXA9UvT9jeszwidigrCcDhOWlTKow0moLe2Xyy5IVYCYIRmU+ly2F
lJ6ZimU3FHbfH+/9x2I343Et+dziS6HYmYelX5IEmHPrw2H3rymxSNwOVsfkJtCJRQBeHQAAq74d
BYDnnA7gCaB0j8YIexxPyrSlMUkhHJAcpBbGzPcqkV92osFdrTgjQsQNEvo1R1InWHIKqoLFrNh5
4XQ0aulaRm8AZnnIiZ4R9gFnZrPyF69+sTRID0g8FA6joO2kvfa2/dAPiG1eLCZDj9VLb9lcsvBc
hKsmYoHCMF5wYsFtdpKI6wLmp0oBvCGI0oW2DG3SDYuK7qKUN3OyA1xAOvmFv1OitfyhOOn4K68W
dxUdXzIhByfH0P3kIEpxgsCsxmvIOaC3I60PYaDED4TpTt09gE7g6LeCZyHNGZ/mYONEwcZhok7V
gklw23v+XHpo08HU5GeCTPn8Jx2CYwyIa7t13DNNpX9NVj0jyuGEK7CMVPwxuxvbbdIVkAu9Yra5
ZnoY5xGAwBszuOkJvrPTcxwwxf/Uh1gIYybH/MEIiR1Yug5t1pA7lORI4eVBRZ6HYPRglkHUNNkR
5Ua6GpYHyWhpVlVxTTOMvwVkoV9FVr2W38IaRHFgJJvhEKIEJrNYg/E4aV+UBHMYlQLbS2fn4UHj
e9S3NP+02AwNjo4POxBUs1pX7Z7XTNmHqX3l7KycNCR1Fht6O8dfF0BunzzctyFvFRFayxfjKnbN
K30SjDCdPH2dpSrSYwToViOcbEoSX2WBokECUwc2I4Fr9u731+Nc6Bv8oimlEb7JOdE6Jc38wY0D
+wlUYyMUxm77op2eLMiZRxHoZvmy4tONOJqg/0iw0DS5rPTOO5uw2WpUfLWpV5cr2PEez/9r75+y
2CmS+W1a+8PsFCtOz/3RbAooib/8WFGj1+0+8nTgYYcUI7gUr2yW0eIC5l+4RK62kNvnTEYfxREr
89AkRw617Wh4RLnyhJY7Q9KsCTA9LHXeDM+LdYp0bdCln2lyF7aXaKrgz9D+F+1Ikm+2EWWmSA1g
io5I9+cRYKui2f9tluwhEDibVZE4cJ+wvYSCYdiIUU3d0HfQKEIK/LCdsEGn0aiJpQPRMa6pSkz6
07jDXo8arnTvqjjM/gtsWMa4uhwdseIENjmDSGz62oOy3HS6mgUu9rHHGENH7UNKGK/Ho8N0waP2
yEUpHhBSISApbM6r7SJyLnHBAACbJIc3ykWqPFhY5ds1k+gYSX061gEvPPQkIqRNXqIg0XMDoYNa
z8jZUW5SeOKGfJszfabTmSRIspvEW76tZjoL4tigmpyCLyMGpu3wNNOHZYjlbomiCo5gaal+EsIB
P5K7G/zefYU0GhGCKOBcQBB2ZNkzTFgBkaUKrKqQVm5aIvamlT+g5rq5GpPkV0OJKYFn5JxfcXOK
G291JJKwA6L+PKHlfxMX2moCJNpS1VEBy0rFzyzZAi5Vc+HrHJeCdcKMhPQRq+MGYUY5qcdXQ5u7
OJvsdi2efgvSV1q8MBUKuvxzHdE3jPK26ri7asWyEbjTW9ZQgrCM9a9mtJ6nuHfkyhekkqBE44jN
Hb1azfmWnovi2lPlxDuDC/tYSIQJuRV3E7V2+zcRhL7Kl/lr9DF8TilsU5EsERrxW2vQpfDGxP/r
oIrmCRXW0LfNl6rM/6T6LLjY0EUZXw0FkAx0IqtPjbuirWnGXT/2QYzT6EYv69FPgkUiGtxm7SN/
SznBQLU7aG+L39CbFYx8H2GgzQnzmv4jf2bt5jHFaci0csu3EW8fyZ2En7CGWO8KJ+WxDIuNucZW
HdDc8fVciz22Gw3iza2jNQ4d4v1+m7tiovX3BeuY4VlLzRzdr8EfKDUFi7KI3dZc8vEKYAn8iDij
CyYV7ndkvisZy5bfIfoZYJEuAfv1iGAcxUioqLTbU3RHJmAU0CY9rA6LAePck3ieECq0iUbbpw2/
Bn3gQ9sZfDIZazJud7WDsH7zGzFSmWNIqDEb2b2cScCnEIF41S4xoIMaDQFAXmIXpvMDLKHbzPJW
SqgorTfDVYx//jbYRk8eIGVBsCCeL+ru+DOda9MXCq2hpgHIHM2jJduBklcfiEX35tKt4fotzInR
KpbUB0uKSh9S6kEagsYhCyzqYDbcecDr/lwrP8LK4uOa6W9xM/1oacp6slNNWPIR4DTf3DH5wX3d
BJzjSRqGkGbzhTWMyB60e5ODZ+0ceL6V4APpB5iPaLKg5nIa1AQxlkSgY/5bsyJdeNqn4tpkDzfh
p1EWM/6V91FViAIA7QaiISARuIWOCBF0DeW8plLChGynZFGjglMAR/xAlUCADKiAW5ashOsxpvT9
DIVVFxJ5cAvZOj7mTfN7OYfavnDT5ZGcSc9eFGZC2npksfOKOe0Ytqiajy/DSZ5uYy62sc3MAonx
WEQE+lGo86dOF2G8JslJtQi5UbcNPiC4O51hVUVBG5//TuJgPB7U02zf9Js7FBnIhPd/HwBBA7TX
R2aO2DPpBXsv/E5eNnXIN11cOxGVfativhS7xpZBJKLLe43N1rdxoyD+vdpQ91ThR63j8WF4l1Wp
p7+bADKRDgO6TQztx7AlxCxsEeD+UEMZF6sdyMRO2acAm2jMZ7QWt/6eXdxCWWmwj+qxXrliEsKx
Nqix3fYufKT9tEhi8J1kNRNG79TyS8ou18RLFdVTO8jMCu7OrAwi9nyWbxiRcimZjB9uwAZevtGd
XmpP+xrAIk3/PrxCW/1USU3Yr+hwrP/1giZ3ijUj81jJkujN/lJp7XLPPEkBHjRWFtgZR3Yy5RKB
pVKDNvs/fxMZuptRgp9bBV64NN49YLTuAx3OYdkRVMGqQ6fTWOkMHf4XfZ/U5YqmUcOsEVjs3r4n
c3jxMzJDzjgfGYOZyWo4w4YuQswDg11hQFfyFKQku/3KUrFqynpo1L+ARDmNYaEZDCPafEGce/QM
g375H/FhNFa0DDoSTG8HsF1JUulCrt9mnYKWHVzyiOA/HShG25zxDY1AwwR0PYIP0mE0Wrl35GOj
+HMIDAJJ0WxGdUDCzNa4WPuYE7LZOOP6VZ5flEZF3vcorAuRLfrMGuejS3fmt0+n6URHY0UEDLCG
R39FO0A95eOYwELOX/YNzVwAKi6B80+3PgJPSDQ35t/NeFD6H5EWmOHCWAuWH0QVxNohpMQVMaxV
ZEj18VQO+biEo4+djPCKDqY4L1rbUfcIGvmBpXvgDcnOI+oJIeDs0Se/kk0jXX8tDH94/RCvyZPZ
6TP6d/VsEJU1MHWORcg3AzSarkaC8avAEoEGjWanPSc3gCW/kpRSoxMdu6biq4wSmJPfgNQ9itAb
4m7KnsifTPTGKv/P7gzLU7u8suXL2lv5ETPYtB6pRB03+DFXQlhwL0RxUOqURr2xVdDWG4bXQ7Mo
6JEJw9mv0UuYIRWpdry8GQwmQWKPF6g0QgdDg4npMyfLMABDhE7QWfuPA/ThkhRiC4gccdfylqxG
jEmHh/YrhpnfryioAslpjEotYhPtDBStEHbsqA9p/H4EilNORoJMfcLaOczw3SpsLfp01vzGZI/t
QHc0vNuipxdSTdIPnxu78rkNavIvJ/kaUn0qPe+lgIZgDAD6REljieungYA7+iqvzLNKgl1dy83p
PGFGCEfwqAAAeuPYUPVmiO9i07PLFO/BeVHSBSVbp5U3eYmFMPapAVeSrtl9vo4KWrH//9NIZkca
T6fmOIheORahHqiAKrjm27TzWxJB8UZJneUojCGgy845UUgaJdKprqigEEmjEqKh5mMDzTIcwOZF
GFXj9RUcWlYUMZRjv4r7HaM/sECC5Wm9H4QsocN8R7euYzk+yd/g6nqyVw7uOa7mIkn1n9GJEHOg
ypjBW0g+rUyPK+0XhPJ7kZjus+AxP9C2OZJRlvCEPknmutTeyrentPcbipb6IanCrT28X+vpfKv/
L5GaJse6xJNz/etrfo2WIGGkjmzerZbYX7KSQP7rH47mJSG8gqoPRyexfGK9cOdYbX3SZF+Dt7Bd
XA029mW9aHlIz8s8Ia1blQ2++dvJujqXlRPWCh0RBCBe3Zq1+qvUtNeDNL4MhG1n8hX3cu9K0HRE
/0Hfn2nzb+dmIjhVIFeUMzLi9V7V0YlTyWihZ/TbK8xVdrtwhAqY7Ly61gXpW+DX/kUde/4S1yBY
JPFbPffQ2Nt4IFlrI34kiZMcqcYR6LMQ3U53gStyqae4rWlijr9R0j0ZtGPx1SEY6X+pNFD0de6X
E6p35UvCRSaQPY1vrHqjVedqSi0czzmG5X92l5TSVh5c9OAoHUd/VW+20jvxwfBB7Le0YFLzR/HB
jqt5kDKJswmX0wu3w/QEziXMhIayubIJ87vaO+oNBJANl3ZhgfB7cygGaUf4lz/JVz2DjGvm2bvO
ruqpSG46ET0KK47LzzSszP7nx5dime87siX6gZ6xKzRN4fpfVWOp6HWqvDdB1x8kF24SCPSUcFwW
zqFXrK8WZ4lQaBcMnh9mHrBp4etddK5VZbkkKBOmvfgac3TXCvN4qjqlf6pIYdg+BUAciwYkCd0J
tUY1sBSEqJ56p+O2qKq93VFtt2pDQtp8p8mP9qTIdKrdnf6Zpy2sJ83vdQFT0rrTUMaXfMMpBIh3
tXuSR4i7pe5Xbn6E5PAeDgULVhkztF50hmMyGKoL8GOiEes++1WhQa0/vSwXCamUl5pJn2LHdVbG
M6vgCqHrkwAdnFBdj9HcRv/4xvZpG4/k/+z2YY+WiteQNMsVYUJjwrloUDpuHXkzIHxLkkhWS9yu
eyLZkjZ+TrE5l8udc0Gqsve0TWH2rlWCNKwimFwKsfy3Om1OQYL8WWVo0eTH8Z30kxpn+v+sxU6M
1GgUCAO+cYJDqDYlPi+b93WlHauBVTLxtO5NBG9/QTBaszktN/8wO2ZQL/b5dr/psBtw6OKiOTdK
Iph0NDMeW1et7j23G7+aR01YQSGPToG+LT3Oy5dz08ZLRNFh4dN6QuDyT3jnMQHy6MJf+OEV4Um6
DUU0v+sCxlLWXFMULBT8LSjn79LRQ3cDUvo6cA4190/BvLMF5FaXlsVcK+Q1ZkDpl11rpQBk1jIj
1yVeRkCoTsdgKafKqs5IC/4145vBdSE+SjAgvUo+P5MMg4jYML5twg2/9kc/3TtWWvXMP17LJscx
XrS8y0/yMfpkcM6oO46FMMdXrxL16FO1g02ymxANaFDv3l29sMoKhWtC4UTPvVTsyuiIrVyaJAMr
Doy9y4MJlVwBqfY1KYewMc71BvVYCOQ9Sem5FdFZPOrRGBqvSxBX8+lp/J9mlJ+xLkeA6RzaHXRY
djmdgORNNbnOm5cgW3peYbjpFjy8FPzaAInWt3bTmLDNFnE899bVmIG+7/i6Ui/yv5u1UnxnytrW
khn1txAeY42GTHAKIQ+Ayfjt/Fj6Ap1U9j+V12+yCfajQZmhR0jMI4znJYqsOsVdaRuRHOpt5JF5
g8vdL99+hVp8EV8ERidGTuvKwfijx3N7Tp2mXw8ozL93kLpKjRALsA/pnoTxpHxXUVgwe05mUVlR
zx4Pz/mddaJc+r+hgi+qtslxBZuM848lUvnlIWmJrsYIuBuro20q+KpzdWQ4ezkEqFIOeopkVl+h
y29HKnBU9J/3uZcfgvJpig2CFd5Jybs05xe43RsqA/KJipOAFlfghA6BwbE9esyncJOarpCTiMCi
kKdzrUYAuIwItFMTpLP+CcOxrb9JYISG5wTvnayQIRVXNX6E8YnLhg0OYcZx862zXjYixfZZX5q2
wCpISJauaXVcUwX5Wr/QAkpDXq8p/EawCAZhtBMEHu1EoPYxzdO0klHPajXlhWhubAOGXIIkRRFq
v8FmeSuKL1dx4Sfm5vaoj/eeG4AOPRsealTDLpVh9BQrk0Xqiuo9SFr0ivx8xDbl5tg2jxPIQgfl
AEe5ZqJJOjALh0XM5g2xH8hy0JkMHq0QE9bClMm3FHY/u6vOHPIwFvQfnpLtJ0pYIKLoYsW7s9wC
ce1QDtuZ4CVLVOk0NRh1oUcDnjXW2tgGLZsgObr7QkHUUkrAm/iZhkIhgzEJIuA5wvklV3LhuXws
WJ3dG5rSyLIGW1IiX70Kvev6HuFNt0lXCz+V3PBnCQdMc3hCh6FmbvDkqM9izx0JqYlDJFAkPldV
81vMDWm2/f/q6cjPtRxA7UV80ZmD0p6dKYk9V812rNdzVMSaCembqWzp/AR2hJ/e64VTk7DVCkV2
RnKzvzbzPICbyRx2f9v6Kl4tovgtZEQguKz/lzh8rgbirV+rvb/Ju7e17Gc35vn3WPpFrdwGwPrK
bLCVv7gmIXnizjVDOMFsL8Fd0IqUyQplTziqZtFIWqGashWuFVw7O574bASrTqEZklZVCGJee4aI
ByVY0eFEs8yfW8x0eGDjkbFL6zBqzPSFHl9cCxWqvAXcxMyrxWtoVd2KiLkOjXZKTk1f96ycSc9b
RicR8xco1jVPOmo9FTqVdMf+OIf1DI0GZgUonzOjs0Gaax6FOVbMGyZ+9+bpmEl8hHFdUvRINioO
LlNU12GAQ7asPdcqBiwOunZZkcktc4ZgrDnJetbrN0yHAzQxCMU00yijnIUvBoe2VycgdkZyKcxL
KkloT8fZS5wS2Y0yb/awV/VFGHd7gklZpM9vnb0o8IejOIfbn4r/xVY9P7WJmk0//uB9/oPdyUUw
7FiK0Z8O+vjN538wDAb9HjKigtuNC2Ne6/KjARRog/ZoSvJsyHz8hoi5q37sKcvFo+fWWzR80va4
DHuxTTnfKqXBvJmmVtMjYRmO45AjIVlaV7N82JDHH+Mc+Kc+ZIMWBuqBW3RxPEmImH0bqIhtHEju
P509nt+6PkUz/wvvTMThlIImZuAWtY498SqM0m24klHzbWVRB/HQUhHC3XOOBd+0mqLGeIclEr3n
f+Q/k3f5C51ya4Pr7RWl0IjOAf8okIOjstG9OxEyb6L5zlHMlchFtQADAJvdB4SQ7lo7hz/YGxr0
VFWhivkv8mDpSLCvJ89PPQ0vH61+thy3ssnnuasTfaKgNalNMQ0SvYQO/2leOxX5bKDJDu5g6kTJ
NEP74KNT4TSvnbwijB6c9S18ADHTdj1oM9iX3+MgrpuBWop/R4XHVZ2cwQKKQ7Z4TUQEKXwT6dWt
2p04Ppk2/DfzfVY87W4QoaNcuXrHy+MJxnNnSZ2QobGPizDechcynrBMPUNNSsK8yiYeZexVQlie
5rft9lHgth3IHQdNTSyZoHll7GHwIyD8leZCZkkuJ/qMFeG/muq+B/l9n93+o7HcQ0cqHzznwQ67
UXIzXkEfZ4QWpHoMi+rRnZMqfgHVe3QyRwKNTED2sp3GVEpQs8qEDf7xY5ElX792q0Yq8NWN2Gx8
nJruvvF40S3AjMJVfQfuqMyedByt8xYK9P4dcD7is9EfM+Wwondjc6YQ7OCJBSIs9efA9O43h/h6
vvnsDcfuxugsevXwIsydtgKiQqu+n53pmZmQvgoqiZSYf6nQ1D4/JHujiSHkreI1zx9ZvNrH/dE+
csFCH3NoLTf6RA/wDDA1oIUN+YynvlPYkciQs6Q15mR8+E/2zyU7wPBU2PaYtG1NSpV2NLQFe6zE
HW82yLlZFhkw1pAvoVfQkEYNvkckL80jee9KrE2zBGU3mN6eIAl9lKbjNigFk3Y+egtuNyuIV+y0
EXImNFPglCA8Sau1LjvkHce5/5gvRHmF1tn21LYX+dqmrFaaezamzcMJBJrdz0roiBKwUOk3qnh2
ChfCWy9NcXsFlSd8kHAG9SUdeBtdZ0VWXjMLkSQ6lW1r4JYX77pqKisN1A2Zx+UFFqUtHQH3k3Gn
qXX/7eau8La4UJP8Ega1h/BxlXpKBl2CkdYmt/R3mNDbvXBZDuGU8T1M+430NazklSEVCNWeNpBJ
LU9sabPpTWfGSDANykMNbp/lZS+/0IB3hSeqXTAU4CLT6q6L+cVZVti6EHCOIJg/WdG0cLwOSI0/
YidaGR93yDyhopumpkIeXihxYmkZtDIhW5qT1/zoxSubDnE+micTw3C9LOU9U9lgFFvpbwkiJvx3
6dEnMWA3HVQuuMATjyJ51v/QxXlBS+TOy0JnYGwBFcMMxwPgGimswAJRM3XCLJRA33+idBFegwxi
UV33arCR5lwpL3hVcaVNDFOoGCLaZ1cI08b3coQUjypOs+JxEuIfN3ASqbYhY22VnbtVtDJ9xwTJ
AucxxLdJ3WZmg4uCEpdygaOAtf1FXQ/QpJr3CEOMmw8c7i9n0mOc5wGwzkHwundBlDiZtoP3iw1k
/lyNMav5gUDKabXgzBI7bKmaiIzQHgli4FF+HenZ7dDoc8LF6Jg8Ws41P4y2ENjJuALGUudPN2qM
4pyOrx0qAx+fLxm5tZj9u/5uJhmnYqf7ht7vjHVLaT/DaZB9KO+AfRbo8Tnrnk9CHdtF/+Nula78
xJNd5Fm/KxHVNLP6n3xU4PPFzhmcoC3CbcnS4xkJ6LTmGyRigRG9YYruN95gTn0E9a+Cslh/hNG0
g13yTlnJOrao5/FPeNsxSrjTI3L6HgwkT4g9FPA9i0MnXY0DnZiXGG+1BToyDlGZBWy099llJhtd
1UQJ1hqZZsNiDinE9jHUJr6YZe6dt6NChC0wXqUipJ0dbX2txqcx5AztN6+iArZIlOp2LInOF1gU
Y6G2sZLxTZZWPs78ZhTTC34vwwJ8//cqBjS+WnqDzBGpikZyeQjq9e7ukxoorL/jZGgcpqqUW3TF
mM6tM1WGG+XopVksEYoRzKTx4jbwRjz0dyMD571E6lnMdPNgGCAoPlrZ+1+qTMDsyjUCfxJ38xJp
/5E8rcztrVwecoS7hrqPd8QQ9m+4uP142AwKzS9tA8WEPtLDiCBv2wMvStVBn1peXoFDN9ODkP/E
R4eX0UPwzTZQUjUhBthGh8eUFDL1psff1ad4Uiu45nPQMZMirxyER47UNLfwAJDGV57PmMh3gz6D
BKTCuydFR1Q5AbHqExR3ti2P256pc/8s+4JYXTAjyCWs6pGLgcikoYH5HpguyHdSid/LDksUEyC4
1OhXnu/TihXS31rZKEs2wXrLGC0lsAdU5VgFZnTOu9CvxPhPtjV4cP7rQsfy7E2lc6+2aj6jE0JR
IJyfGY82SP29w8yzIiLRGFOKdZnuPZx5jn0FWNxGnaUcO4/XWUCyopcScqEsWPJInsI7+yUD6/Dj
GdV1nTgyjtnXcNCTRW2Ln9ppZMwbIPIBItrHOT8Wb8//Gft9VY8fq0HlotNWYwoTlQkaHh+q89v9
PHKndaibdUnIIcC9rtm8Q4hvrCNirQLBZS8RiRU2mpCM4mUBtJJRwz17UpLL6IvEfHqcsMj96Kkg
kzpuffUihJeUJ6Whz/mbiiBHp2lnJLo33xH4fwP5u763DEisDL5avswH7sizbgpm1omVio0HucrR
z0u1Vomsw9TYcK/fT+yMlG5zDRGZG/nH31JsAlHPJRF9lsfBgGF/EdSkTXjaTweGeFZTl+T9x0gK
8OyCnZziPz/cJ2tixn0YAF3PntBQVrsqtiyP9wjFSgFX/tO8vOIBdib6vLIEY4Tn2umD/BGV/yX9
zEvdJNH50PFWkp2ECu2fzTjYxJHyFB1s+7fqk54xcQWTyjlIrBRATM45xQRM4hqXvI5eMwlciCER
SdAS6QJBTJIa/rcpDkv+2bFfhVXT88nMic42SokvIjd7BspUouPsM7TN4oHR8jtPOMWF3f2jouRR
E0NBmZ1MzXQchbZfHkUvnDb5342WvYxro7qM1wuemFVJDWZM10QtESjT+Cr2egiL142zCemW9dCb
ejEewe2NoP+h0f0iQiB0I+XjvxQ+oQRqoz3IGrRkwxBBlZfjguoMZHYoaDSNFuEmrDBZbrISNLy/
fv93RrNciZhekLqTVF14z5czEmx9KM1gCnYcDFY1CLsxtTmNNQgS9hn5Za2ik2yQbBvHgTGaJ8RN
SUO8mBX/bovYQDUwffjvx1Ju8Ou0PA2mZgB9+cvMeLzAu/sZZ5C7IzOoBTurmAKpp+ZjkAacVVCA
0AscUdtZcCCspIm3pJv4CR+hQCa7hqK7ps5fLICc3uo+HyiDZWSW2hJKCkQ7PQ3sg79H1AjGsobO
1jR3LudafAp/IkeqrElHhAZOn8BJZse/OrQqZokIF6MOne6OjJ4NwwvHpcEk2omPIWZoX8QxYehb
A/LZgvCRkJ5fV+PUeWEMm3Dq+iPFNQJiYhq+Ai4GPbCo2bqSMpf+YB5OtFyiIs2UFL+hcqETGvQE
1mgcFwH7mOSy2dRTbaKEDWKZrKJ2JU5BKZcaUXDsQOBDN1jXTqg9Vn4SaM1OqIh3+osAyV1L7ziv
nWMsbU3ZSWnESZz44UdMzSRxIr5+uK5/le8UoohyrBF4QbVTb9iYTAC742ExfvGDyLFlk34hvrdp
bsgnOBMhhnrN2raLCyNiw5QV8FxSMaqAxTKEThoqQ0NMtL7zogERj+rVAc22uVHsrK1tS/BHoOzz
NQ4x4vToU3KDXtKw4aWIP6aA+MUI41KbBmuEcqBwpAOyMIXaCZsEDxjnKL43y/QvNt8KbdrNFMQg
IuyjHpSXHcm1BNJcjrwj0Ou1p9F3nvJtbnxKfW/ljoeRt04uy9+xBvS0Z22N3rCpN+t++4D7mHtR
eA28T9bWkKA8tgkSIxtFyDpAORIha5QiKOKJx8L9ZO7sN8enTLKFsDwAyoiqYnD2taiKAyInbfBT
i2MJUCFcYoM7IJZgrJIzGJp6/Jz2pty70X2RYn3g8AAWPiNy7b9QOwnDX6UBpze+7K2A8vNZggVV
VhI7uKRPZGvfqOZLYadeqthMJxNQNmQp0O0OGMLFjR15gaWz4cu9U5GsYtBPZaARs511+8w+YYP3
uNNorNlMAYgdrqJm0fwsqOhKhPTdrqTxZ2bq1l7s6xLJ4lP+TeruB3u7KP2gcdDi8S8kh1PS1xO2
dXgaTsrsoG2112fn6fD7pr88JQd4Zn9lg9O5as3jcIBtX6A/TUxPdmjqYzUGM1mfOF+dyil8qVfx
L9YLQzNz+/36l4eFa2l1egZ1tW7O4Ep+AWnd7yCwf1T3mWYKM4rJjfQeQIXpZKzCJsnw1xb8o8nX
AxuIpk25aD9aBcKnHgFBkFluV1/7opAgYtNa+jHFyRueYrT9jU4o20YcFNLuQj1N75qoc/kTFJxy
kEv4lJ7xWJ1DyjpUK/GOnyNZXdTfylqS2ABA3VMKsQ+oPT7gbQ0y0H23zmyW2PsywBfuntklbh0k
PIkcQlYaTeLwcvgLwHh0c6x7iyuSbB+KT72wgKnKsXavChvrWDz4+6BeQ6vxfRhyCKSRa/B3c0bE
Aayad6MPg1AeIBe5K9KHFLlCJWWUfPDpvZuDXn0EhusZbmHQh1uOWM0YVq7JagTJqofOLcDOGYSn
CBzO2VvLXLtO+pszgGBuYXrVc7dkjGHa9Z2MVyLHo27hySJ52q3wKN4mbQqmvuFq9yjD6Vxu5YwM
B4/mgZSgcD+Hs7VC1eXc5Fy6GRAujmSI3CIv0cKvA2xoDLJ13jyYY+E8QgtAIJMMnr/xDtoOA11f
go61vCHjhWsDrpjR1W9Zhlee9VwAlN+U8uT/jyazSJ042xEcjS0BTOuMxtUFFMOvRTbD3tPOBc/7
LSvh5wdYq76mo+wao9H6XxLZL/WMpvxhXzw9Fz7C31fkji/XNnlhxuHh2LnMmgF9epmZ1FHPOsTc
aT+tbpk+OxF3bGZrdzNUi2uGFuGXuV094y4m4SCvXOtoP2y7zgI3BLDQQDZVP4t5S/I5NxLSyPQ8
C4H1nYVS8sqyXJuFBHpUzlO0LzwpNbvXpyjXBRmCt8ztYCb4mEs+M5wnFuvNWF/UkgIGAdI12Vl6
j6PSi3eygQgtor5t9Ungj7k6UQZZTlcb8vJAMeINLUFBhQJ0GvTN5LDxFC2NlnvhEebRUuinEzx8
fg9lq7aULHBaExOAJSw4yuLhd3fGUUUsjiJcSIwNJdTv11kYhsuP5F/kAhUemhaYnlkhosFp5PvC
p/mRJtBBAiSqYctzK3Ar24sfXcll9O5KkAPxtpf76TBPobJkntxSHvzTMHwwsuZuAeCxKI4W2lbG
QEjUcqCuWPCttVlzgmQ+iYm+cxGdmu+o7BqV885Lv3P8nRZEayavG7la2DVvuQbF1rCbm25NUXyq
Pn9+VK3h+zt9bb4BJ1ywGKs/aufIzVdB8yN/PyZjxeJTTlKsxmxBt8Hnl+X0qF5bqtk3TlR52tsC
sKSn71MFP+14ONRUfI9LpfmNveCPsOCihXD6qDm0+5GRWV9xwppTcBcXYzUyWxpsmNVJ31p4N5VO
vPESI0fzRaSh965wtEs5WcT87TOJlbjQnf5JXiFDcDr8OfbhzPQOxl4jXkzDcZBdm3eKwJKVTzg8
cD6ssDgSy234kuNy/QTApsBwoV6+ve0rfv8oGWQkynFtNpby8QHjyCpWJ03e9R/wZF8PHllskxOe
ppP5HSZBPvapyUadq9ZSweVKlONy58N6YUkdbrLJic0dZ1Xop+cUWV5kYHn9i46keO5oektnYx4b
o/eriEyoCvL1tx3NBkdNO5bl2taWQVfLpL2MvD5WfNRMXTHUfqLWHhtokuoXhXNO3wLDCNnXqaFg
zptpiv305F4WnD0733ZvCAVR4bb9QjmNcgO+HTXnJ1UyDX9yBgUvXhPwuWJJRCwliCfhs8CZapaP
YG4NuJmsxncfaOOzmT4jyA3BBvdf+A9XMJ73HiZ5s99sgWT7P5ysKMk4nJAo8XXy94umlHguOGt7
Y3tm/ral2OOQ2SdpZC38NRLx6Br+lhMS4idH8jiIQE5MCVZeiSzNURfEHWTfttysaV6V8AlcVlMi
ttfiA1C/ppvYiUcXYxN/94iGSneVtlb/xkcebzsoUq2NlE6WjLd1usMg0c/uYtGMNuZIBwEtMjMY
Od07xOgAuVut3TWKJSTTUX6zRPN3A/z4wWK0RQM6clOkPlJn0qsx6r1PU1ctijH7dk2Zp0OZrxwH
VGaVGXGA7gQ6H702uUBt0NE6YWnMGKvi73mhP/Zz6fI98VVsmj8aYisas8hDBv4s7YLfyN9tNsMC
u8DavlNBrZsDpqkgUkJBrsr+g1LyVFgeTFPxHVqp21ln7FYg/TIDcLp5jifD3hCA2wrTCzSpOUIp
ubmwpIfFoqAWeSiVLMl66p9wx6AfUGWVbjGRcfHKRUrYm6b4CSYBwpUBmIt8eYlyMh4wWpkacboV
qAAjSgu4beOvGKrMCPop1DcJRf2eI0O223/wuhBZCgLXOw9i77Thr62VfSFEIqOimhyZ5Y93cab0
f/8m0t0j7UZ35vTWwJrq0mZ7iYJdxVtuDYCfRxiSt+R0fmB+/1UzOGNGWjq9SkJbxB1JhSFDfMrC
tj/c2HpV48YUaL4f3XAnD6fpcDfo5pQnTTmwABY2p+DzBcUp0fmve8pD94eFe0Vsu4kFNiI5dnu1
8CYlF2BGTgzOQCxzRQzWEDYY99ixf5yZ/IYAF1zRVwtZL4kJfdpisc1H3caHZLrWm0jJnaDOdT70
Nxugp4v1TyRNmhg1Nc1OkwY9R8S2cp3Ecm3A0/NVYwDAIFhJdmdRmJU+6B2JYJ/nFQfMBBl5Qod4
GzR8nEVwNiUZhX7JDbH5c8iG1dx/5UWhC9tOyX0MspYyE11tvXTfVo7nOGcfg1A9KsYWoukxxkrN
aLl+guBRCf3bgBGK+F5i7py0IVq2P2/cU5aUzp7R+wJEjTx1tzyQrxI1xa7WH9nb6jFJdZNUmsc4
Z10q+Vb8r+ecK6FMfErmPrBrTZR1a2l2wL3AVX//FHF1lG7tj3ARQ9gGEckEtg6GSa3dNJIoFSWR
tJ/KZ/QNSEs5dfa2rtQZKgTwp9mO3jlIOGX6OnRMIbI9knG73AeOUsjknneX4VdVzU3jBTPMDjMj
N8ywnBn/epEXj2cvcCDFO1sF57MG6acZ8JbK0Ky/7BZ5oR247D8TpQtwfF5pKlQbQQnV2mLrDWyD
AtLf8zcwnAcE1w1KGFZgVrX2vOs68r4Q++ZP2Tk7oBbxYlNL6829w0SHfjJlK/JQQIBUszbVdR9+
7+7Mc8r/G+ssrBtNgKj3UfhxKci0lmEkhQu+4Pe2yucP8rNQZZiufjUH8MlWjYO4xsQX6P/0uqZZ
7s5VpXwAO1ZC48yJDFbatMxDdN3S5Faod8Pu1ePgBj0Bi/hdJ6/ZxyYEnNwf2IbHWYwYet2sy8p7
bDjV2NY6y6HgsUiAPJ1wnovuuaPLB/KJZZqspatCUZt2BVB4uP44cE5Wrw/KrKjK6Fh29+jPZqVp
qGyeAV+cIWu/x9bgteFs6cw1y0H69YoyxFyH419U/SMqapcNn5hlM2ET+8tZ4oX1TNQV15ehBig2
Ocw5HbfvRkpC5zjNLcsDcfEiSo1i8CENfhhRyuXwFgfntYXjsody3xB73EEiq6RyxtqSyh3DCauo
uMc4waki5WV5pMFMsUC9xMqQVWoptSsXjUmrrUYkEHGp0h1Ox1TeBcVhhcSKZxeXiCvtwLP164Kt
42G7PGWXAEWu/ZIqrHHdFG/8GYfIgZcOpAG6kiBtV9Z8uVPIqen7V5R6uSW/QX0/JIAv9nQC0OkJ
nmUzjN+3rXjQVnaHN+IZzrrF4kh9Ut4ydmEbwWyai9gpUeKYfLvfk6wzFGp2pzdSfXwta5asDBpL
Of/mt7IaXE2VhEjlKuDvAS5LesRu0EMjoVRy+jn2X+UZTwdWY1SgAvozx6VMdB1mZLcEc0hsA/8O
YHnwDlksFEM9QhnnV6b9RdgNERart4dgsMLVNL5SaGghJVCzAYMJL5k1DWF53iOOjpM9XIM4wjMX
5PfMybbJD3TsQ8E1AzRrbdj1V3AMUGvMykiFYFIDtGMx/gsCDJ5o5eR5kmxi59HQjg5ssImilTny
PQenS3FDvjZvzSw70SpdBbcBSubA3yQaIyBGJPXMVSWGBVlVAhm/awYpfPi1RQbGKkSsDazX7uqe
+yKROPjSZVpW6Jf6+IjpFNBg2cPlsi9F8lPeoyaqFo58mT3K3+2gi2EvRd7KeCcEiub7lIeTe/gZ
BRmXTMmzoh2cZxoqOJEY7gvfk8D1GAcX0mzHE3v3ZKshRMm5cvOereUNKTrgfBchAhblnzStB6W2
p2HmttaVV5s1d7SuNz/L7vOgdr+OQ2rnfLZv3cHcAfrYcAF9hMT7qlwBk280jctqszz5NX88YvGS
rCGvMkxLQrNlvQGhHTDjd3LXKAfctziB1Jne7L+AROa0tcua3/atkeA7O42cnvsd/bjZjEHxq+si
uxWtWFWGJnRaKezG2A9DfDsboQ4GlLak6mOhnZzuJTe68mGwSX88fHpBac+vZXWStwyCJolQBFZ6
1xWwZuCzwKc61v1hPzRXnyJWPSqLM+6KU+QIuWulF/CZW+9ab6lpYbmb04Fv6aNbH+8wSO8RuxKf
kJhk+TDhuSWzRefboyZS6sZ3C8qq3IVmj4pbpq5n4Yed9bluhelYdRE9lNBz0S/4JV1VoassMVps
jc3eSbPvIJqN3o3JwpMwEtqvjQYysVxJPYOwLPaojD43ApEw35qu6AOJXSyBh/0wkfrGr8PCuTjS
q3grM30+HjKEcxiYevYzlFrWQdLqs6AYmc+sHn0wTifFmB/IBm8i8qZTSoJ8H7gTxh6H9Osl79Dy
JhCyOiTsLKB1geSpxvnM0OrHiFwBbyO0W72twWBvuv7hrCxznPpjMZ3YuRY+7J+IieYaXEkADxc4
8JYf+bdj8Hft6F1X6RIp34617odPbA3KNOo22huCtsbSxh19mkPKHu6uhY6wOriEZea0UA27fS2o
4sF8eBeSONDYaTaLKgqK26g27rVjVQdQJkdi+l1r46TQYi1azmf2y6mypo1ANFVudNdYm4Zbd83e
nBD+oQvoz0pemRw8qZxnu1fRyXDTknLTY2Oczw38mrH/fRFlU9B9njn3PndEaLM2KKIucCeV0R8v
oi4jVvnEeWtFQ6UVUyakeCLXGihN8AtyaK0Lcvb+Mi3xONjOsmuEeO3mR5k4Bru9kavdJpIH1MfV
Luocp8Kvpkp6zZiVhUrct2lo1gZkjI5k4L5PZ4umGH/oExJZ3PW7O3gwy/EtPTUCgdt+S/vJFhLy
cvNk8vGse9BSWh68+RzSZJWCr+4lO9uMl2OUNDZkiZlEes6Y6wXRgy6wT1SSStML7vdhjbC35HWn
J0qxi7BVpaxMTe95R1mQ8OTr4xGGwwmHMw4iKOSZ8O88LL9WezVmw6XOdCNCtDrcIEvMQ7EsyWS2
HaOK636fdd2r6Ki8tWGQCcKVfUI9ISUTNKdgkblmENqZ8CJWha+zynvUY/REkBcDPJ3dVxG6m9ku
VHO+BVLdzH7//j7d0j+CbIlHBf+diLsl8tlhYevG4yxA1ysmGsB/Fflsaqk8V3iGigSpVi2LG0pO
8dMkO+DWATtMpSzDvThty7+BCtdvHUViC4Y4BZYdLyVrwaZnH7GIxn8LO7o67O8WO/qRnNnfcO02
O6fG9AwuwgpzQV4Xt89S+Gul3JnGd6djbQQhK32iuTs2HKy8r/g8TeSJiABeZTEDTvFtnUgS7L4G
zhbevzpILLAAC9yahzeWLAxnmoUwt+WAVtIzpa3OeqxtHlw+kmcV2FttFmXuzDru10OON2g4H2hW
BYthpxp75Cqg6gcAO/yrjoV5rYsBXj51R+J9AibpxFO/i7xqpCEQ8PPsOE6Bn6P8T4KvVxt1AAqI
0nPluqAbwCHhO4D1mk0Y9GyVLqWoOvuhYzYmpRU4i+RbCpCe5KNGa8TabAGfLCueXfQubqMYLsy8
tdwmQudZF/zd15vezTfi1CmLKWxZw0os85Nx0vBPWZ04cvo6I3u/nwiXBLF2ti7XUplpeIanVJmV
bNB2MHc0ZI2Kw1IamPK6U5NOKua/X79/81Lt0TO7/uTiVQpKy4WGa6/TBh3olKIU3cnZPAZTLL1C
ZZyK5FJKxLcuMnicf9d9afq9OmjyFlIidW73b5E32rmav418zcBx6RNe5xJGS7yq+udhL+vWLSPc
eXR/WZJ0v5IbS/rPh+BHuueLMn5BoFnbWIFArmlveCV8hF/Z2LdoGmnETpRm+xjU21/HVD0Hm7b7
BRO6J3t+DkA5NvOxmrIoPcHY6UpDbETqv0AQHTrRooqf+TKdfiQApM2d0jh4JEtKI8goyOhcWozu
dbd2NMBP+7jzPI5bECmc/dBnl4+5mVnkP+hKla3pXAXstiOIFjBHBWsb3LNNWyPxOqHKeUfd+IBz
r0/R+VsBVouPI73VdJleJK7U+0stOb4j8fLLY6P7oqYtxmJ8pMa2fY3paioNbDRzYroa/CprFswU
0msowLmxcJs7CT7QTgagkphcDFWkyri5DFl4PdHhLp4xKhT8QLkoCwHkv3AL2fi2vvuqPx4cXT+4
N3Yfy7VAsLPt8G+oiQg7Tr6LU7hOWGERHyc0c+r8hacne5lNNQcfQjU8KFK7UR+oC/dmHXpDhhj0
rgH+Fneyhh5VQx8Of7CTbPuJTQin065uBTxjkJ0B55vPdOUejbWWsbgVqS4u4qh92u0VIHU8Mhyw
q9qkcHetWr4pprB65WAXEsa17WtU9o5t9wmYbNbEhU6JPhLFFQBqiRDujeraEIVjSju/V+FyciHk
f0FmW7q/bD6gz0Zq+QC4m3IjKDmvpijsEb4IB5QHAyjbMOFjsF0LVxJYVS7AIyKxzzZBAXJitk08
n3b5hahfRjMoa4b6wtdo6BE4K3l7xMhDSRbG8/7PlHOKVrIU08dpXXGRYNTzeX4UCStc/RVMJwV7
rPzGutO567WtYayBd61nQpshHiEBy8y55Z78VdwM2pfJi8I7eHMmuEIi/6yRbqwAm2JjMZCVgpTJ
wX6LmLD5S8Oaa63qdRgq0RAFh0FtQ7wPNa6BtQRuU6nShyvEsOEdvhrTxCzMZqX+RzSeg/kwOnbl
Fwpov8RSW7A+rIiOdCP7bjMkCWNPoxubmqrBk9OIlgzV5NTTL9Ttrmhk51IRUH58B6ptoboimtgm
Q1DLaIydzWtZ8uhLjlYOAp8bxT04dw1Ake12Ir2C/XtqUyRnF1zoZN4Qd2kgoEXmotl9DKRk/DL9
vYMp4y9MxxmLthdaErOzuzwpsW1fVdO7ElQD7eLpef5rC3TuTS+1Zaer7hlUlrD/WHPh+xfGDXub
Pvfeq0IJZwVoG1XsY2WLyd5kqCk221IXIqwA6+X/nwNwPx8JUJoA3/2Q4v1ydH+PkDl7r9IEfgu6
BJqPH3dGGtNZkyrMiB1HVM4dmzZlwGailrC2BKPTcAvajzNWLoovPf/48AHbprBerEARtmrD90ZA
OUh+rDKqGZXYgAgvLZXrmLolgH7W97UB5iuggK4Dh/G+eJm0gDiNEnDXgouH41GslAww6TXWPdk0
unRMqIiHIdcHX8PJCVkVjHZqBuyPAkmyKS5YUXcJKbwjcDyVKhIIiCrj6AQ5DtLUr9RV2HiofZOP
Ncww8oC7IAxP3e10cbnqqCBjr9RGU2LVsX4sD6zbUfcB0IoDjTVnCwgkceZ5Gda1j/gWjWBsEOS3
TNCdxxCSY7MYBEShAvnM64XsZGrcUuvHO0VxdOWtfLHIAoAVHMslf0sUcgyCoQktD2cV14NWNHx1
05l/Jzbsto4duc2FdFLyHy2xcGLsEJGXMKtGM3OLeGJEthdJAZDDdtdw0lehtsHVu9unE5xIeULt
NPGFf2NSygL1i/cei+LaL/4OGhD5dmffIq6DJWWgxYD6mMUQJJP3ftERkMJF6yEqVxZnaRvB+aLH
u2E0R1gkjqtxwod7s7Oo08OaldDbJQus2Lu6IMxXBVGDGJWyaxpGphRAg1zNAJqRgdCqArN4wMGe
/v1FL6P+WH0TBJfSFo6eORYIGuDHQUJ9bJY29gsZfd+ZsDYBrITe8NWXIId2rhYMoLFsHesQWs+c
c4VYA6MmcDyKpINsGzPsDNdFSC5p/QRIOR1eGaZZix/QWe6NT+oCUKYTwaDXsM58hnoi4hNXgyll
0i+ZGEJW2AYchUrf7YFCVvkfJrMR62sYbjYeG6i96Rp4uR67E6JNGrmrAm1Y6HLRRaBP84LfHmcY
4Kb1Dz5NnJlD3VcfWcQLSdn0t21eVfIFMKncq57Mrh3IgIwdBLSfcNI+8yt0GZZbscxOzahF5D0N
CgtS56wfaidqIvI1/UE3k7JITaP8rYLmazzDyuSZ0hj6vC6mWs/Dm7Od/dPnmKseHHuYcMQjg+iG
Ag+yQ6v9mxiRj2hjPES+ZZzY/D0R654kjYiEohxXA6yJDn/7gaaOZWYG77oySVzfscf+SxLd7dxz
UT0J7OmfM9fxfKr7MkfTSuH32cCHwnf+OgTJferi19vFYcDlkyB81tS1MMekzxFzYPr2t0CT75j5
OCF28+5WCJQiDL1nuijkUVlcYhfiRf4Ih/MMbreHW+aZQ1MVHYhb4B1iajlLnPRf1YYiVEzUBe4Z
fqL4KwwvxYwt+KJbTCEZcG4xC8a4pHvYvWe/bQ6P/wsAhRgWbhqWAjwujErDWmpWZOp7TYmmRJfd
qDsn/Nzv987Ej2zufvuzjCiPUloyNwrpkogcO3PXWM/JAKz3/1+43oAhHLMAbYG6NGOwtipYpyy0
GkloICqNvr+uKv8QT2pRcoqf4cfgSjTeuUVLf1gQ2oLfdy3UpQ8i/haJC12WLMnFHFZ79zz6UNwj
rTmf3voHCTChaa716cO90n+G/MTHvn7QQGQ3jJocWu9qBFxr99432bOF00jvbIf8mrf9Gy6un0li
PzEDLaufaYz0qsAMC7A7OtaNGVyPEAD5BFHtbuHH4olcR+JnfdcyVByvyCRlRXdmCbvyEjrtUqRg
s2SM5+iFaKYh/mw2ocP4lP977Xe3sklNZVPi/MXZFNWiS7B8hJ7+QalzWnFhAgARBrA+H4EIY1FN
SIugKY8gi7FVSG0k9l0ApIS7En7JNp5iuY4Kz9cbwWMp3HvhkDRvKlM4GYWXYUp9+1856chInF9C
cSastgmIbvH2JT8Rb5rTG6ilRjmLGPAFom0E38X+OdRHfF6kY/RGYoLpUL4rUbox0A6WbetDL8Ho
i1QfL1OSlyPkdtHgWo+utiKxEbUtB1yZ2jTj0OVZH86K/lkOsrbqogqEDYtLb5P6tF9YgvU2Yjfm
/3ZBS8d/ixzxt/jkce4stOd+BPkafFUHAyjOjQCVhsHEBYONxc2EWJioYZ5uKDjkaLhVKo5mz0FG
A18KCj1MsoyXyGpOz8h+ioiABWs6xVb6yp8KBZ+sMNMWFwHzOPqKW9K0wsVCHow0jpZ9PboxU76a
jS+6JByos0yaQHFivlqsjv/oXet4sQeydT5LdWRTNVr7LNAy7gRA9F7nef+G19vBzgAPMk8jbVb7
DTa+LFnVPGOegtLiyFxB3T6zf0PMLBn/2+c93QIU98NZ0hDt2z93105aLTP7asbL80CGEIlXc7h3
O3x7ssx0k9HF4Pc2J4JnF2ov+NlANiT/gcGI7PlKkA66J8a8SpNp7Wg0FvqOMKgmBCxTtvxsAZV6
++y1akeqOChf57y8WJ7afe/5wQbj/1xqKbfxcs0MIBobCiJmZXI+kJ6kJUGd6eGobYPOy8/MR123
kNMQ4elG1bjgib73JIOLCnqkRH2kyqalpWahGUZn2teUX6HGb2ZDEJHssUe3iZmVgkM+6GXz7/af
yK4JqA+mNIQ658RIYdcx0bUUxKAnIgHzKUTmYonAECWgriNOWnBdFuNIIx9kDIt8D7m+vTXxPJMq
iS2ZN52SV+Xn9M290ANq9GkXMKA5xLMsN0bbVLkaVKx/gn7y+ivaZtdFYgYUg8ExNqMPRV+ymImR
i9I96CC2rg3Nfukrs/8bI+XFI8+7eKB57gBMTbpwfSssdo1OOBztp9wILtoQyPGnQ64iVXafusZo
H7jeNc6Dqgcbe10QYqLgYtBkMxxVpL2AvOEPsmW0cHqwpYqCkdk0vbg5bpxGlL2itUcIQndFQo+S
g1ot1shIXS9vvKTpY557SuJ3R8GhB3LThtPp7S4XkDLjsGgmnTiUPXt1mr9US5y/+kaC3Elm6Rd4
2ECGeBsw4SEMbhMzuq/A6+y12LeS1yIws8vcFYqoUxPNB9LSI7+maF1dTXtP1UGwyMkc0f7DnXK0
Szbcur00Cm2tzarrmbBwYqmsouLPksSdbj6G1V1GaEMe2XIzWRTku9AHbRMyBFmMnLJAwrubv9UE
hTYl9Ys0DdvZgp09H4aOXpD3t5wNe92LYqiEbrKadv2DVixvT/NLQOLwHikxQnwQRY6pxZm5IfkA
iDOi/pkxK2waD50XOne5WqnWBkEvsvhKcYs5sZSbblLmASMKREReILUOJLqO0uIneCvvkeS8tC6u
ytQutbiHGltYjgk2ffvnLR+kRIHYDgmMxyNidLgddFA8v8ccMkSQiW/NhXsdL2J+SgatHrtQACpr
q1uX3Mii42mmBNvm2sYnGOzgzOGCpKWNtNdTGPNr6O55PjnOvH2H6KMhAmF4U0axx4qlExZSJ9N+
dwzKCMnJazijh9sYaIEs2j2fPVFT6HYY6mMONPEh2aJPJdo00zlxmpovnPKJTdo/cd4BxY6m2SRo
N6bzTkaK5UQxV6FF+whSODQ+qlMtgceAqZ27o1eT6xb1LmmN3xCtXrRVJmQBubb1ZOY77BX8js0x
jYb50Jxil2l7zkdj8jG96x8wRnGGHRXnp9NFvhBf5ACQac9T0PYU/nCNsbomBHepVyJNlHOHE9Ug
VHfQz3vqXszhUC0QUn4PuCxCuwqxUBPKgMLrJE/LQocHz5zM0MH9AwH3JazsW0Bl/Z4XYRvUY8BX
UzkfoUMFln38eUY47W7SnhxF/eedGye7yC0//3IfyphwtdG9ghUhauka21eoysY7UoGlybA8mcP2
7s+OTstbI4oa+54zPl73Q25jrv4eG4srkJuGBpNX31nE4YnofTG9VWcc/ekbyGOYKyTHxiMZ9OmH
haRxeNlJ1W2jjlYA2IfhFPvPM+9TdaIkQcoP31sgjk3GG3XHEU9aU8JpRU2MbNJ4BqmXY3DH9v8R
lbkb+VHc1yJ4E5VfQ8Fdx7eEPEVxnXqR4yjodLVUlpSL7bOAbtEvaJq3BvxcnkHENh13yii8ocJ/
cFSS9pcooOr/AOJCpTMbjQwqI+OKqA4vH1MklHvdmvyW/Un/okpG/vHFhMiUKuhsHE2XyyZD+Kn5
JvknPbCV2T4ZJSbZNPFsfngotff3q3mrAYCr85E8BZSa4DW4W6i24fJ+OevFDNgjO69Sl8l1yVBz
FUnqAoVLLEdQKUXHgy3GVlSXfo9tTezhZHgYYv/5ETBWzX2aau05ZfS6DXO/fg4KffFv9Cj/1aNx
Dkezs6FIHlMOEl2h+52X99BIy2wibuKxtUOeU4rK/xe5H7+QPhJE8oePjAgGgwO6/nO3hwOTgTcX
jdlksXB00ARd0crAGpSY8k7O5olO8BbVIDgmYSPE/D1e8ZKKqmNGAzbzcipnCBRHi7vxWJwd1bcH
4CVwPLEB90IAiG/RNXytxZTHF1d4Jw2ymtNBFvMYoG0i6blyyeiakWjw649TAjzOphmzOJTC349g
zxeiAf0Fdbn9SuXOJc6DIwgh2oRDpObvrwQXFnf5Rw5TUNDdOIXc8twHFTxjPrzKGpRnYL3UyIED
prwXl+Gt4qJkNxe3NFfsbBAkZjbCPQC93fKFONaBkvJ1FNiEj0OKtoha6smvRYiZ6bQWhuB1xtjW
oofpqh548CEurw1N52PVI+be6DlbeI4TAgHRYrj2GGELPqZ6XEU03ThGfX8hTIOeCiL4+cLZtTYt
9F/7fcZFAnzybDQainire2owzo0X27aJeWMoxo7OVcb6+ONWHCfJzfWcQvwxl6uURSj3JaFZC3CM
hhpPAYxtBLECMb/YVJ9ZLhgp6fxavYgRIj82lOoL+ns6Z2WBZRZKScETSYyGT7IK6T1mAPqywlch
rsFXun5A6lz533SN+lUIdgtB6zaJ4buvjOMGC7v88Ef1R+yHbEkuwHi7Mb+fF4UPQ/aW7+REyzzn
WwCOCxSFKWFjZdVldpRacNa5AgFu17+Akl/GzGeYaDJSpPstHSlm8d87y7xEpPm/mZ8pSE/Ewz2E
X1ooHXxMAu+LEFamp9WBcZ85JewUlH1kYjcfEggrOKjAP+KFHmTsgzp5jZN92y+RMMPe6RhF+KEP
dK0sg+Hr9H+5JEAnvqRO1HvA/UAlidnR3Fy8RY2brTMP3FWAkxOf/LfMT2ERnUbkI6OQPlkBdIwW
RaC1My+b++DkN+kuUdB+7QxPzvpGJkT/FIybYHVL9SyhZqjL9C4XMRuwhOD52MvCaoN5ZAJopLKR
utVq+QNKzClVZx57B4pyUSwovfYfFQmLFFe04fUq0Yl2P/xhJkPgnUWRGp9HWv1St/1zJPpiOKUR
DDi552ZCub/E7aOSJ8v8XrNQcPW8RhFKvvZ0S7KCF6U2hEb38rdjRjG7l/8IWq0Xz8mM7XIxgTsP
kn7rf532kfde6KP3N6ogEWR6a6iu1fG854akphflI+3WqsmwWo9NDk42TGTJw5zHw7z5s6eEzcgQ
GcX7DZ4DuLiuAKZdEOyc+tRyVmPf+dB3EJMSxEUZHraOXHFu6BeqRHxayjsCDsIiL9h1WErTzWgX
KClCHCy3NIDe32OEpEG9sfHvVwrF31Q3W9S1Z9ufi4JGD1i7dtA6bIjVXfyXi7SwaOoN4ltAnuQw
DPHYjto1ho3Nxc7aYeW+3iuMHtQsD8ZYEkfcZkREODw+Xn/S7b9JA1KqfuGKQR67q2GgattLJhz3
gLphc1IaWtxa9V2PR458d9uP9gyi4qbKTOPO2pYTlXhhbtQn4n3ap8Bil+BRehJR/7dkNPXKewAV
K4HVu14FL4Zz/zNNJvoj1BbosHJudlN9tSWT4BfU8SBsYcr2AliYqGfwvgDH8wblNSTc5ngv9z+c
BGFgUnee8ucaoH9LzNBy9aSX2M8WlKA97mgV4/z5aiBNZxwo6Kp/OpKaAg61ioBGgiOikgRhty/W
rZTkRZyFSwQtFb0iBu28dmrhTECG5lvzwHfDC3arkG+dPXsm/oZd1nyzO1wbQZ2AW15GjmAm50tN
FfmWGlzhEaq/78jMV6YIYNkHx8JVZz13vwpPTK6dC3jBQmlxBoXYO5Ud1FcqByrxE6YigHo+/y1s
up3+Ea+0Dbe8hCwPHYFMV/Lgmvkwzt6TIxWNEoKDXmbU1v7KZni2uD/g2d7sFdapwutwvZ8/tSDN
35wD4oHIvpwGC88WGTBCjFhkCQd34EYRU2VHU+4c6XTK21r70qrSOfjyOR28GBdJyyjn7/X2EFJj
yk7fGtYjVG9iS94R5B/3WI+xsDEL+E7Ct2iw9E1TQk5m8IQZnUUqR9pinE1gUTdv26/si2H2uKKl
EFjigmTJOwz2+jT83Yq8FnuEP7GxDAi+aMugLdHAh7k5ems1nbukxU6LV7JtJ6BILjKpjJPUOOk3
PDugY7i+eB1YklfBQH3sHwA1jIC0nzN8Yy3YeVQTYfubGdln8xmjhBiHEL6KOAMjQOryNDbRvGrg
n7E9ZH/IS772+3HvsycDqLByEb5KXqCFSf+dtKMh2BQKnqC1LrLKK7N0H4aKuWq8B1RcapnzYcZV
8+ldDaglhaCSPAIkPn+GLohIbu7vYkLCpfwfSXwVxIEh/Y73Uxf+vU9QaIq9n9xQjSrLh1O9nxdm
GqnytkJAFua3f61uHWvZ/twt9qp2mrYIfxSPi16qHcLIq6oObVQ+jDMKhJhH2THzGzLVa40T3i+G
LYYA/yPQGJiB335/s1wjEr3vFiaJAvQt5IIFMFntASZZPVObZfJmE1637jyk9REMWH9EX2J2TcxS
58MiNc+3FxXBaEw5ZTQXymcQyvUbRXurWRSToa+61oremf0cYDJwEOSUGElF5O20dB81cmzRvNAV
D957pKzIezVqQzc2+omvdcLBrZf4p8OjC4bFDBKi0RCmesn4Aj4PDTH+WyoMEXkavw2Bzn1a21dz
eltMe9OQo25/HBQ7HSHuNudXaCMzZrrKghA5Ueguzjc4KEeAzKcbeHnjUtzYQ6QtO++Ox0Hnd5h3
Qo4B0MXoOGTJ+5w6oElYE7ugl9T3Ken1p+5CUtVhRc9pn16+fhhITbQKWIeXNpt7NKoYFFux71Cr
kZSH1Welei6TKhqEhPfQkfYD8xmhjTN5x79tTv2zzZ0+2R4U9p/kO7+JDfuiCg5feqnGUcvK/w/k
BGCzGDITbQKBNal9VF0NMy5Pdb8fvF0a4H1Dd0X9PaTWLmOWwX5iPcHjYyc6DjMNkExI9vkEKdlb
zXHx3YxXimkgrF0GsVMSQe6BDhR1ROmeEL6O31B92miBqLRdogkYwJyF/b13pKl9TfRcBBbqXzOX
BUAkUEF6v9cyaMUwVyKtPpEKG/TIl56th+evMXnPLJD28RswdwYblSz0hk+VNqYWhsBoaZr7jka5
Y65vliEyD1Xj7nlZD7u/Rc0lAXlI5Bwc+RxcAMbgEl6rVYi6YtQYil1L3DQdl8TEOlH5Lj8glS2U
F8kVrXgPxvH4p5wWR+LgTfFOXDArWDagb54+f9lFTINPhYQOi2MzBFEILKpAsqm0u36ojMzei3+r
vkbx0oeNyHzRyM9z3/RHJj9mF5JRPfClkqEtzpqs1us+3yKDlYdqeAx+N+tlIFAnGLjfaXjJ8YLf
eOegMElnozZ+2CJHIcJrlP/K0jj6bjMVBQ50YdPbAgmwU8oLx8Nl7kOVebJwg2mrmy9b++BhSYHx
MEj4rDuAbaBTa3RFR9XZivvBQjALMCrxrb/+WLt+dGJ1MikaZNbj8bLZxoYFIpFQiYeENFdxJ6OU
NwAXcaELFU8rjp3bz7+KZ2+4M0VTXJ6rut6HZXgpXqUdlHmmJOetx/qXshIsTiju9dv48CqqJ/pW
Hm5KHjncLESYLaJnxQYXIryUrmRzHgXNG4gn9aotLpckHv+JIV+tc3yqBAr+1hTZNNN9dMCiaY7p
Shwuni9yjLOp72UjiGCq3c2yBXbYeTnhIc4iSXDs0KVLw7McpVv7zQ61RgQjyupTGDbzsmpXEVTh
201xxZIHmWErIBTyB6QrCdcV1bXrgcoLhFYXZ33e/jDGmhOrRb5YFdQiZAcoDouP2IRD+FALubpx
BBbzPOSWFqmvXRt3gMaYc8KK+apelxN7dUcYwPl0iuM3PzwQ5KP9ZjzsE6yWYXVbrc/0KYytzQbi
P1J7PqlZl+6FvWUqL02lj35Gz0lMeMsil6q4B5pbLMfACxSmgRcjODmEMoMaCVEk42sbUiUgO1D+
m2a3OlyCgyJKNkGcDoLCI38zIX/52Sid1Nv+fCvNPUCst+AuzmlgvXnadxiDJ3t3JylfhpJfDvM+
LsH6jpx1I6SmJlrrbLvhlNVdiCl/JuvYG25eAtyKqbgXnBW7coeji4SfOUtegfR4QDqQYngCrTF6
eByqtmwEtcHKAiRftf7Z067Dzk6Iheu+U+hk3wj8wxn2sxgbxThiYfnNnZ/NrRZjXqzRj0a2fI4t
KChDvWUGNbAPIUoG9n1zCCh9/6fti3V7H0aeB4x0gRQtt8vbzj0eimmPpEdWfZokfgh5j2OKk7p/
QHGRPkG2IxrsfLxAP46Dj7iZBawCnBcYhk48eNUvFOz2aCsuOhiW/ozdCgK3o1g0e4A7XlVR0y4h
yb9xBYD/CZY/Si9THOuBOUUocdBmv771UIQeZ7TmiC/eSpCTTh0EtbE5/A9l2d0RGUy5/zbsl+ct
FXbyxNM4P+i7lU+0XyaLltim2eUJuRZ1hbxmIHoUImbqiV4xb01dBIvNnOz1tl5ALEI2jHFScb6r
VR/hljW6p5mHhb6gCnTDVnGqVToXz+RYHnd7kg4K0xZHZ9FUzD1xi7YpZ6id9c4uaU/oAp7Iggq6
l87sp/WbfidRUvQd4t7xJa11YK1GFEumLzyJwVdtkHKZqoAH9f/r2Nas4nIGNz6/h7fL4yXXCrDD
GbWyEZSM/+wvcVVm8FESqr0DQUR2v4gzWaAhCUDMPuwASeSvZDS9aIfj09DyVVy8Qh0u7DORIMEp
CfHpeBa3p6zqbX1eFT1HVqeerAXh9Hqh9qiyJhF+Z9Up+QkXrgK5m9/0yFOAgB1ZAGsNfbn2hBT6
yYdC3oJK+zm7KCY10Y6CN9+yEBvj5gbmNoglth1BJ7nTsHte4SyXPaVOQcAwNgQnY/3UEcTO+MOS
7M5dMWxhzmMwLSiMlZ92dq7IoiNJc+VzwGJwlcVzNpahiXcS3ZnP6YnEiI84jHGU9eahkwytVxcC
grxCYWNLp47E2qFgVwqzGPtaqP2pdL0FEEDufWdX13wotQRSvb/1NigGYAFUixh/kyorIWbf/CQC
wxy1jacnCndLl5Z78dT6oU3kQi0bErQutQP7XmuWJoMyIWcCtGix20grUGLk9HKj0pBAXoljE912
oVNXKtg4r2Rdec/EyorrXF8tuWAqaeQ8OX4CrQYIrz64Zz5JacivPBNqW9SM+fpQ1chn5gr0NyH+
uvjy+FIwIvlbaKxGVxKl0aVWUjIuoLXldOFiSjE79yzhQaoIUbHZ08zIwmBrDun3xoM6Dclqoifo
AvGjMpA0jLfas72UCeNofWn6BA8Kmd5Qc6mtOZYpGPC2Zh4NrHBp2jvJkLsmbWQK/BgeBOw2jX0O
tMu1GndwCt1V1vNEQcSb65mLMFPFPEed2FtLbnXSkV+ufwEx5Xy3yqZjIQSP8f20nplNKDpZ4G1R
DGk8qdXggwaqQGl44SKxqcqW9OuLQrxxemja4cE4v7KCmhD5M753veryvDFk3d+NAv5QId4h3lEJ
ztrm7gYLXZ4W15NLw+XDK/o8PHSK3KU9MLJ6irzLU4oJqsY4HinKvqSl6/gFzN40jGb/ZtIJRJH5
fjtK+Vmk1JrRVsPlsYUVBKwENAvnuyTvSV6Hgls5trzhDfOsMjI9PxvwzhbdWJddDYmTeYkRCz4Q
NIf6e41QBH8PjYf9s7ree4DNXFMDGtFJBkbwKc2euF0WNTq8e1oZG2eUvaVaTzku+bTlQhFx62+c
QA/9RgoYmjs71vEzP+Epxay+cUTBsyrqyncA65XBkJ937SlGLJHr9MAN16XXf5wZnthghVMgV8/P
Cd7+D2hKzsh7/xBVmmqW/iA57d2cWavz0ddxWj+i+Y9MEeiSY8a72UDSmorQLg2OnOc9A6EDP2xi
WYImGSHjP7NxfQ7Raf+xpuQ/ZUE34L+BIHEVERSvYSGU3w3S6CYYRd58ABO6EQ61I8egQjr3vwv9
JD+bAcCX4Jo0Y2lfDUPCtAPdMaeEreVBQQXqfGJUHDYQb278wxGS4lPfgnxJ3s6Wx8GTI26F7k3F
/rVJvZPp+kCM/WoY2a8OEgD8mwCxRAFjx5saYotcbk5lJ4J4uXbSPoxrgnff06E95y4HOSlkMt3Y
gAlgXt2s1kjwJ/zYIWGscqVRppugBefNj55f6RqHttaWAZ0HhX9fdDxnG7fdcmAiPRyXuDA5xLZX
rxNjeuMtllp1oz1F20UWcezPdgl2GimzY8xoFagfYHKeKVPmQFURS4AQANXnixLtPuXWJHGox0CQ
1Ik0A3/LeCnm4b1ZAr5v9ndjzP7YGVXm1ZljTd0IDFIzzxRhmJsk3yqdJRF3Xwurx+LxZfe8BRII
Lc5+8YC5sGqFZUysmZbNTobYqL+YtUZQnOcTkwdCwfM1vO8mXEe2VGk4mb5RVtoA0yWzCrsKEFKZ
j6RgbLMOv7cNNS7V2sBYcUJjVm5Ww+0yaDdHs0z4/pEYQ5L+hicdTJT6HiMiLmV3N92CxhMudBur
2pG++X1rGwPXXbBtN3GeqQ8kK79biCUUpSZqZVx7igtAjP7BO1sJMqEQfxE1eyR4IhVVyx0HpaGN
UDGiMcAlXbTOIW6D4bqPvVGfPNF3K6T+9Kh57k1Pqkue3NXVYbxE8zlGgroFv/mi6pZWHonJtSzx
5mdhC3lQrxLRNwGPsMq7eKecWAlO3ltflDH8ajBpUgzOYw83yNUi0yp3MPOaSoYbSRDsnCMhI2kl
np3cjZ2g3lyhGePhlIQ3vYemQ5JhJUr6Bgfy2QKBQzdmJ9ZYKl3oErfkEuLXYuG12/V6YvS1SKPt
MrW37C8cpAnyeBalcI4evnMq+Q+A6J2IGLdcT1BsGpw7OEVA1EmCo5EFCwu0qg9Jc8IB9Iu8qwPg
KLogavyP4oyzvhKhrHfbdTjWl6NqFMH3CEPMeanZ8NUnmq8Upg3yR/D7rMwJd4mAMIiDA0+v2QXH
PFtfzvZK4FfgW+zQmfZdhJyjZ9H5RUMK3djQid85pe62jl4d9ZqPb8up423L+V/uxOZX3+1Tfd+M
HtPugIpeC1wbteUG9u4bkv6jQb2qi/QXJRC1fYhnkaYVmINrNXb4oH/fgCXTt5ajSc41G6qxKDe2
hSVOMgmjTiYseTJF5QCNmkrQrO8YQ12bJiMs4aQQ57RVLOb2CfpM/npyew4w8zj1PMuXLHakAcYt
9ebx+wYDsfNphmL97nallUbQhEAPLRMXjYCvuSwacRf3brF2ypugZ8xkqlxVUtAJZwM2fdV+YQcA
ANgx+jTNep+TZA2vxfYKbcbZhU5WMLuftmebWgyrfNghwZTioC/xkfLcy8wyEeL6CHH0jm4vZOMN
Ju3v9vpjfxAbOOK2VAUjbvx4CY1wvs60quLx39mSMAS8BfVtvALJXTfT2cuIjczD98CJRII9+V8a
JLtev0ImrVlgjj5wxiMpPNJzKf6Oy8CbmMHiMYvdZkU0nEO1kwPmFKPq/86Yz6j5C5STXjRroFBw
hAGVyWptqrm+Bdq8wfgu1uXDsFObzPijSIjeo2pHen6ZPGA9CB8ziUgojk8RPcndxCinQzyaapAN
cbZc3sDF4rEHb4Vc1mqF1jd7WSrRFrGavDVND4F17RkaeXORo3IpabtMtmxqlm1quFeKCiUByJsc
DuyD9eFtpAQZ7acNOkOP9+DjMiC1a70b3KoQog5POrJVsOcCNX7u8Rm08VE32u0E1ZFH0J7BBmfH
ChJ8el4vZ8vVdZV6PoBcdjQHINpV6MMSSmKWVMDytWDDndKJwhOQykm2ymNmqTwzaiE8nzcLP6Xj
UiuhaosH8UUoVyFIH8FBnyiVGgwpgY58hF8vOhnANZjHLyDXtGrYaXhd73LLIVjL4HzkowgwPxAm
ge7CvF2qrAivJjyi1AB3c2tJA9x2CWym28q/gkzM0dHIHH/DC640+/HVFweAp518XYeiPDgGBMGO
vTf9OsJYjhmVQRUcs1lkCR/rKSwRsVcVDe/6lS0PpzG1CVavkAo1qWjtm0wnp7rQ0p9kxfTPOgT3
q5U6dDd3CCf2GtN5k9VqiCfm9Dvw1Ph2Jq8clpwiuEblQa+7H6JskgCwCHtBGAIgA62uK6vkFlt6
cTf7aOCaxDr+RPjm/blY5OuHrixBku0Dr0rx5P7CvgPtPhSk5yAj42GB4D1QSwn4AsoJtRpoIpnZ
XVsKj76XPBwMJUsZoStjVGpl7JJhQJCzT50x708yi31gB236O25XpZv3ygAbGzc+Y9hnSbv883vh
/pnoz/OsK2MDqb/NMalQgAC0hpZgx1VR+UWE21mb8zYboCFgMXg2r9JguoKo2TWU+YlLAJvSfVHE
yE6LjK8qzh45YAu9bn+VSyeXKoxLNGJvw8wSPDXwOP/IuoKUhQ25pZzhp+OX7v+hyA+yP1xTOJzu
CXdUjlvU4tLTsCzfUlV7gVF27oqjn2M8FRyQJsyc0vPT5OEQ3auNTnpwpmNThYun8H8rLDnK4XOw
2w9TfcA7FMYnG8asGwRC3dWXoW9gGTvxZBl6V+07pSYdNZ/1ATv2NVSdkJWMTzw6sOa3io60GD4U
3wdT3jIRKM6iWY/jud/R6gBAOsgLF+aFD3XBljCMKhjocNXsOK3FmjNCY7g9YgA/Kh0YOdJ9gvor
9ndJHgTkQVMH53clwYfeZAwxFDqRcElrXbqqznSH4cGum8VmC+zs7ZQjOBOr+cuJe3T/EMIShG7o
9Nm4mD1uMkQgzPGAQpH4r/5wDp/mJwc/vjXAoPBFGpUlH4SYzARJ+d52DAvxPGGtvLVn/8PTvPUe
SzfgJ3UrglqBZUEpkB/pg/VB1YKw1Em/zoNjJcbponFXzvexTRMSlfcRWMvPIpiSpXdW7aJLvYxT
TuawGBwe7sNgqguWlQzvG2B+m7fM4XLru6I7jP355Q5QLK0WKSxcWH5vMqe7rOhAo4Sn+JeuOhKp
R/r7L/3VmSr7wqg8l8XuQHzlzMQvVa5jB2qcBT7W/TZDke36OFErDI35WXYlQGfrcMKkB7ttnnMT
KUtYECKrylezbreLhB+ZpYbIYHM8VTx0A6qba576GvRpGoSiZYHXSoFKTMxJ4kEn66UOq1gVwx8w
3DEwNS8bFESpWI8zeKFQ9OxwpYqFFNRYTkr2+1e9gVziKjDld010pnq23I8OoWuOcrAnljt9ETfm
glMZYn5qBaTaTKFsFRQ0lrOYySdbJAn7lYy+sc4Bj3DuFuX/DHGB2YasuVW9G8QnbHsEBTkAB5kt
m9ZxtuZ1g2wP60u1c0G2udlphpnasbx7ApZnOq/ZnxM29YQNHRnNVhiiMylDpCfLs/nPBmuYFbZK
Q+qvbgr1m7fLqss5WDfiE8PO1SBbNmoSlMPjKS2rtRN800HTfFD7seyktFKYpDlmBNYcrIdm0gYP
JY3XlEXGFGgnUBgzths1Nz2VP3D8G8H3MyDfjI1Tfkw0B1NFSsvWL2ZJD/3z/QHRK2w6q3LjbFNm
qUNM/wsEORnAYj4XxbOyELQQNiFMdYsEWsHNTt44MxYdi5aMrD4RJY3QfZezZrq67BbbmU+/U/lu
YQp42SUJIbOkmhy/SqBEL8xfxS3G3LqRy4rNMwJNEMziLlis8HhU5Hx8IOKdQf5tUqUpUfqCHFad
TMDnzHbzQzylhAacOR4r8d0T2nNeuYp6XreicjdNTjkv1HGSxeTH8nmZrE0uGSNKgGRlTXh4l/YD
LW/oSlReVQTZZ/j52Wdw1cH9hEz5DmruwOoQ58Cv06wiPaPcKD1/qelOoYQVHdb9/nj8NYNqQqxY
rCFdoyknQJzqqIdhIgWoY40hgdWtp4amNA55tZkm067EPHa3vXVN27VGgzK5YEPN+qj1xE0dMzFa
SvRH8ovDlEtS5sDJ6gbNGiFQ1ocrb2uVfEl853xfAgHmwGgik4y2FFDr0BDPf7U2qaCvQIe9H+wz
sljYdhSgSaVMgGLOfJ5i9NFzQaIp9w4IuZH5q9ho1WxBGazaimhiKl4lmwTcuWaP8yrieT5o2zg0
t1RFEefm3zLornPfQqgcvBFAMEIm3XyAj/3sOotKreULvHs2l38Vmg5kwxNVupsfWKmmF4H9WnTA
P8INvCKk87Hp7YlZ9BFXWzTB5pJacNa599jClw9dAETp54h9bzYHtln5aShuYQzcB8xAaA751Rjr
NYmSwdMAuron9laPnVPXABVTQ/aXD5sVFJiMdbTABLEC8O02Tow3RwktzAC3zdJKxhR2orcAxxtq
upI5a6A3FPz4JhXny4atB+7DJdypSmB+4kXSQVWlvSP4667JOakkE+FN9+WTjhxv4Ad3XyeEFc6i
rjakJ4aI4RJRKUgDjcur8IDiHAsvDndgvyAUkeQ6UrXVtDXRLtFpHjwqLr6XGULS+stwgNTcnGX6
lvaeaPj1gLTA0CJkq0RVqbUAtEOd9KFtQhzPyxDgWAndlWuDVRSwTZODpwFvjmw3qykp4ac51FBx
d2bTH68sDpQ/o0vQ+qINXJEnLHZpcFQsG6VkX2XlbHn8HTHVTLuhsmhQCcQPKqaI90RFhvc0VgAU
vivNIqt86oM6YgoP1tv6C0gYctqf98oagzmFONk6pSDyrOGz7lIuhhwfBcPoDRwcof/nR/O4fCL5
+AUF4H1IjJbSdnqknN5vpS1uySSyA8Y0aBORdarxuX+VD6cNS+vh/uN/7aCJzFts5mGWbhALhHa5
oGcInhTtQT+vQc9G0a0ot1s1I6S8tumJ7zhONYFcZYYFU8o2YzgM6zcgVrxOUNORzAp1XT3bXFP4
XL62yodbqbktmXCPvYYeP+RqZ70GiJt7qGc9skM4OI5uYlMB1R0Dis2uw0P94lKOtQ4lWjL0oEh2
Qta9Wp/3b1br4ozcjXxuuXbLazp+Z3FsFK8b5rzCAz/puUeZZYF4O15yewvBDt5yOwZldJ2N6Nce
zgQhNX1fMGMlqlDmpLPcSc3wNAU22tLZ6whsaZzLTWvAwo2EKS1g2mCc+I3E6UBxMzHwFnhrhkH1
j6LJSDTpvkpZPVy33jqmRZT1mwtq78+EtDGgKv95pakMRzls9mIHLSMIgz0BASONIsDt7T4SC5VW
abVtPO0ClDCDWmcOsiiB3oeDkZDtzdfiG9ye40QkHZpy27x2sZiL4xA5rrUrbrXLYDyJbl2E/Po/
ZbMIwt0MKDo1GNoUQBMVVIs4ET3V94R3oLFb9TLINdrq9yBxNa8O8ux8Y9Uo5Cm2HiRt92KIqCE6
kj4M4cXqTsned/uA6QCDvZRxtoc8krN+Z9gn5g8VDxfPdgOit7UT9HVcGDAyErDDdDX5D/qOWfY2
O2IvOX6OF/S7r6RRcsBSTRtyq34M8xetpZAe/6NVwiZG5/zmFz+rFLMJbOCok+OqhQHbokBUSIje
R7KhSo9l/6gbmq+ZX85pZNRDjrIsUzueUZoQkYprD81r7NN9a7EZG01aMx+zg1sIHYkNOVhutL1I
Yna1khGl28oItITi/ptprDt61xicbwZ7c8rg9Im68Cxbvwu0XTErdfTFd8b4Bt4s6tgpApb9nJ+O
W/VY4f3JRnbW129pC95v+O38AmLnw7n6hziZCE1/uum+e0tatCcX9IxMXaAOpy+pv0Aq/Qaj/L4P
M8oyoXynhn2tlUW2P8OXG+mAfETjRXIpDzacVv1UAvbORK/RhXGgUJ2O/fW6MNgQRvOE+3/t5EWL
sEsDmwVvvvEzPcpEQA2oXf8yJINCU5DsOe0PD3un1zFFU3mdjkfuvfXLLng+KkmQYroILAzEcdYL
ir+np7mrqpXvpRkC/XNMWQ3xrvOYaiu8vxLkTLq/9/fZzDinpAY4o239oJuGjVWJwWLqyrj3xUZi
SdjWzDA/yb64GPvScOLAQOq0DntRvHGuiKQOc5m3q5Efo7ZcNhLYhtLTiQEBVymM4NPVv903EOO8
VuBGV+OnqamaI2PD446YbnVdGWf4yMYOKriVoXBOJUhQMzFpYuPr60lkWw+pxuQpmxLbqR4KHZh4
IoRMUr0MbhYkQvuPKlYUIR/UiaIZW5v3dXtNTuC2FJSwLjDW9NrHDOwQByGJIYzjfxcmDJax+B2C
ha/dipgFjVzVBbk8cV0pSBpAKyedvRsR0Yc+4Vd5BjTDm7F3yPI+r2fy5NBF8lK+XUkucGRqoRi+
atUN+7W0JomZlIbAAlP5QKJsZlL56oW0cfdkIweg3d+qmbbf2HvJ+rqW9QP41bJyLpRfWy0OViPu
+Zg/kHzA88HoQgFGk2qQeMIefKdJbpjqz0V4bQSxRInv98zWuEtWtAxW9DmGfFtlcjDy8AIv9C1Z
UV2xAGdyUDG3eu85N+rNtY012tgdgKpObHLYQYSEBsR/Ea+2Cmzm9kzcxWb6XzmuZgzY2nVCC8LU
ulfgyhYi5XsPNnOl9BtVuuunHz5nV8NRolsFlxs4IwGuFZbhfch6knSFW24WzVrmiRcj7uIVBpJM
IJF4Zsg/wheBcUCBoMgaV1y8Y59gR+tV3IVG3wloYwiJFHmCeHxXrxTbm4M5x+q61ZSeElvBZfMS
5AdezFR8qfzOsNdhoZDJ0sA6N0Cxa8jZV7fZK+aX+2x3bre1PBjrZJdUbVPZ7lYoU+lErpOPq/UI
6Wl3eghWmPwNG+FOQ+5ZDchpQVWmR6JzMB7vqta/9pF2Z/nwYm/5MzciXuBYy/Pz4XwV7Ve6JO53
sXAzKy7MGwHNMuDD2FWb0Zz9rbDRyBMHyoAk80hY7nimYIOFhnWfP6pHKi9N0y751VQDfqnVurJI
bE5CRnqF61S8iM6DZsvV37qGrOTIZu4Gu6FN+00NKw6q9jRbkmMGmSlYQYIPuJEA3N2JAkf/ZeMO
mib0NN78Nn5L5DKI5z8a45xVBTFT6tNHkP1kNTqCUpJ85rizHfk+NQMJv1snmSxffG3ts2HuUEmv
wUh8ucmGYt1K/2gAcfHxMy9sBHa3l/OsxCbLRmmMGxWdtl8Ed8IFTAGVRJHc/5L9XuV1eORyUiNW
d/J1wkprnSDUJHDTTOaSR2G9mqTA8t55eAE5T+H5O3iGM1XMSjQ5tbAIvFwIJv03kZmZp8fOGJON
7VlvCZGbZg++efTVi5FQ/uhDz6CfN9vjHmccoxE8zBFPlZ0OR9gGuDdt6j/P14Bo7ERs98N0qgvp
dupYxhRyk5ijsU55r/biUDTeHrNuO4j0zwmrP5JnzafjdlD9kkYt1dRGjBmL56GXAz58Y1B6Ne10
2FXXnV3X65YslS+rrXw2N+xCk76hnHFlnWKT44GxoxYCKMJ1x+a/NnqD3V+6sK38s4XAH1Mj2HsR
uQkrdBgia3b+VnPu+es5DTulo82YVkF3qE3ZAde1xmRXZGyoosFF+dje2csUdJ2pj+Rt0R4HuNX9
2LRjB/esjQW/jFr4Wb2ntvT6E87nCCzBMbrs6XtiHlgfOQxCgMnRkiMYxx1qiJH15JPCGf5POt05
mkRNAAJ8mo/JOq6zzsfBVICtoGqe5koTE5bWwCviiVe/XmY9cSKm31bDTfe6hkriY50wPzfWrdNL
HwyO033dc7eM3Uunp2/bOFBQ/+nSGV+/vHRE5bkFTME18+tmNhHNxUeKMK8xn4vLKEGgR3aRCh+O
KPOTiJuch1mMED/0f8PABIzCMC/B4T0MR0x0iJZBvP1EJ9YUcBn40EKGoMoKA0Q3IZ/O8IhU2PN1
QHbuZbHA2Jn2wQBx57AKwrUp5fqUeVDc0Y9qn5nf16O6TdWdz1JL+zKMNgfRgVVkUQ0vvCkFjlDC
Zv/pPlIYnpGEBlV/SVWuGWyCoqKF+sVEnRE7vMuhDMBsoKHMChDzPsD7tgFc9lQTh5znCk/caYLr
azwO5Fo0CQCGa6w+/SDi4bmTPNblyRcEZAbhHW7VwGCI6CVTfcCT2TH+8f9kQ63HXIuYPNyTre2l
8Wcb30D/runagFuHdCxjsU56IRJzGNThmv9h2Aos5WpL7R2QAOjsKGn3dl0tIFTEY9TvMq0lKpvA
xGMuKKOJgwAj+89YPcrpFhOZakvYJi3ADCX7sxYjea1wHXNnZcyTzjb5rugLfZHJ0rVZCCveDpfS
lUMsuhbh2c4O4t333Y6O7vx8iLHCrd/pANWAS06vIG2TOPtlrK8LqOwbrNtv7s12csgOIN5f18+4
OLtFE0VlLGajnxLlmLEsogE4AyIlkuiBtNnS81CGZxpVwwH+15cMxeI9fjqNyeIrb2Nu2+03iv9V
5X/lN9xAtUKv3D/HGpvN85ucA6SVUWAuvBzp2A00GevTTC6ngSjPIU07krGzvsOu6ehoOR4FBpDg
GvAzSLVxqRa3lDEiwQhGR03DpGL7UPpyk9JoIKWCcLifzqDYH/uscIwPgs1suP7lDArWWcotjFxR
y00VhfR7aFtOSTR9kbyBRJ03nxxvxdk3EYgSPV0A0cAF84kNFiQf8neXjp3gP9ZJk+i2z9Ja8EuM
5BbhjvzKKeQQjl0i0m6yPvjKZD4T7dmJUZVzRDJ6obo3zHCCJsD974VTDZuwsrsJSueFs6bQvpjD
arl+syQ570SUqnohNtuKVDdOUXG8RspifQ8R/7OFbttvELDBm9spQ+9maAE3E3GKGjWNsRnJoQQx
s095ZsLg5xBDhke5NI3DX/AM989CHYF5z971fONhKv9Jy52MtZiwmpMou13b10BLIMcdk9OZSZ+1
V1OKuYWfy+HtUT6jhRTCRvuueOIiMb3FwVI7RQnJy7RODH4neB9JTdEH5t8Y5YAUabuiQz4LM27s
Yseaw2PRhDkBvSM9561irj0wida+VTeuIvaUpgA0Oh+DIe67tDehFc1rSehTTm5Oi/0PL5t2VEEI
1084KNz8JFXkB7JF5N1SvpwN170XRBlvgpjVBwUuNCCG0wu1H/Q1mP1f2sKv07msSrMxWcrQ15f9
1dzEVGGxHxYwedOczVWEC8ljmaQO0DeT7wui3Z8MBr63lbbPlVQg9qVbT39cqcUtiNR3Hue+darl
82Fh1BjmO+8Tr7rkBT1n7PluEjJB59+CJP8Sc931Xc3ioUSlaDiHvelKG8NrZf5rjQBNxHLqB0Bq
gDVXAQJgzIe8KVD3NMuo14TNiP28jXwq3QjJkeXXci7+HwNzBBlOij8WYLYvD7LKPKa3CUn56WHb
M+udQlPHj2MmUOmtsIZ7z8SG5NjzQ/X6/PepVSbU1b/TaAZ0IlW9LFyC/FHD1zo0WnOol8lwemgh
xKN+hbvyxQnzxId/h+UD79enzV53ECm46G8jkR+Tp3PqNZoJEmT0mkkolz6e4/2qjizpcoFp7dWr
HENsGaA7LRiqGUPzvy2hcoJOYU6KXRA8nCj/xvomf90rpx/uBKCB7zxi7utU+EYZZSMlPEYLdfPV
m698kabjeaFNoip1huMXH6YTiu21d6f0iKORH2V/QGMzkcuQCectoIs6+RuV1VomGE5HWH5YFiz1
iDGITNPn8b/ljCV6o+wA2TOpsXPiK1V8+5omzX/rejG8VXN4w98gkZEtmzTx5Iv4/JzlPaDdQiYN
yT85M17d7AQ5bXQhicbsBdTLk/K+aI1npQHRROU1Cym7wHQi017VwciIEdENEYEMoBsdGZySgrQX
P2XeUBnf0vaiW/J9ahj35SMi96SP4UiV6BzBwAaMkC30DpQlaPGgTkj4yBgzRO1QPCNKls2hKS+V
yc3PrcH/R7EUxreCLAM6jJ3YUoQt62zW2w+EQVzqR2mAfdjookFm04WCmZRCx76zYQXqYOUcNCDB
q4pblmcJU0mmtVQeDJCVuhzOf+bY1U8YkUn/cLSiSMzK0KQ1zbSzUiqf7cTt7aUO46qkfD1eVYkT
Fh2yvSxL/Xmf9sV2p8gWoxwA1QMRDyjLbtYEpthw9RejRe2jdRodTwpJOeMeBtzaiGvA82DnEOL0
6MkkQ1O6E9NXItpC5X/EDH2pvQ5cNAVtvVpdgxXdwn//rj5KgXW+jkMnA/6MAeWjAEUrBdLc7aTX
a6VTka9TgHwQ3jdikByhsZ5RppOf8vikesrxL4s10ZnIZxeEkRBIGSjJVVM2rw/5vFKMVqLUjxX5
DaacdG0aHkQm5rWgKpDcr6QnZird7Buesp80hvWLORv2GGqmBUId6KoLeVytE/NB6mwsE7pyevOs
rqGr5e49xBS59klrBGLZvT9gax8IMn8/uR4LS5b6ruTzvDBJEeV13faJtMGavTIjV0moY9hN18V6
T7RmpF6Lnbzh7w7p33fGzsb537Ci7EcBRzJeXGPRaBQNrIaFXJX2P15CuEK9dBRG87yrVeyUqMfP
q6lsmZGYz+tXQRnMlkVrEXKrLg7MF6KVerWEOMwrIIaAxXiiXs7ZxiXuj4dBIIsIpMxe/z78WA/X
/pu2GRM8AGQAUjnTponkQZNkBlE/EpZ7t+K+wpPSF7NNHEAAcsls7Y4jJdRsHWY2fyvcouGnkJis
OZc8SGO3Rd8OROE9+yVRcc2QIc5qeD2CbM13/SemSm9vimlB+pQ/d0uwpyGJYwTIxGnAhQGh80Rp
4SeaikieCxMvbe0+fsu8DOYpojw+UInCsUesum8iMk4bvTw1qSzIpS67jGqiN605OSB6KS9gqYSt
x0e4kZJiHQC4tywHpwkJDwtXjlr9vPma43FJHH5UrsMlYqUwKWeSPVCEx8XWxPiSAQAazyQoFRNd
gLLpwyzv7FHvrdMbQpMj6gsJ1XIlOSyLPu8RO7YZ7wAFeKE9QwpkgT/g+XhGNXCibOF6dN6d4LIO
wEmx77bLP7GUdhzoS2HmHEHrMjuh7Y1PdmWocy7JqAZHI+zojKQ8FVklb2rfWvuJri1tiORrPOXG
SmGsVpqbXt9FhwYeijvsOmAUgj89AIHXVY2uNAf+7DkMshKY9CTnSPKiDDQ6zFKbeWjJzR/OYfKP
82Rtw1o0IR0Cu847f6sPUdNkqWUWCUwpknb2zsJXkEqPn6b0SPL/LDP0BIFJY//T6C+N4EfI5ZMa
a9tjkwQ1nda0N6zKZDKy8nYeQVu1yz1yWP+OqCOoK+jbxj3FjDDIDScWhTFdy8eznxPVIIstz7hp
zZ6ETZLWjhqnUOwhqBdfKC4k0WSktqr+34fGwY63yG8JrHAeaQHyWjf5+K72PPqlrDdAdL78gWTb
lEinZhH5SkxwGN5NlYIJ562GlD0PjsPAQMWom4S36JVOJ+gLbOIkCifB+q/pwcPVJH8hOYaU0cV8
KV6FMWI2+d2OKmbztvNamZO4fL2dMg02rE+cpRT+NKUaVyj0T3P4rVX0gAemsVLCY6EwtCX55EPC
50Df0YaTzuOHQIC0dEjXNXrMN1VhxGK1o00NKVIJ8a66BR6nZ6XqVThsRbJIwoGeCgMgl6SkZPwX
nFbpXC2OuBoR7SVAAghtN0B+YWUD5MDjJqMEcpzgc1hI0q9GV6MC/ldSX+Vpj1dffoC71eoC0LJm
FrrBUsAqkCXPgwkZMhPBJAcsdjmlvBaQMlBsbgYKCOAtcep8Wcic9wN8xXT6caRM7mH7np0Bh6eM
tdi2xWeaqdx3PGjbSS7m3bejc/zDynXBAkIDN/6bNieBCfseJU+9vV70ZaQwrx7dAAIdNtSwYdSB
/1MBU+c6HHtPMYsbvV/VbQ8IU2g/rDAdy6Mo30vqky+lmT8dYyeTzPaqOpmklkiqjSHnfuLmG+QO
oc2PXYdMwa1cg9qV4hHRdywCGSNHqrSBwgJK10vEdnkwM+lY/3ujANe07JSslHT8DmmXIUXlMLQ/
I8mOHxQsOvBNamsfcnACbGs9CYtTl8JOjCU69YxlHjQD9g+XCB8XyPHPYod8iUpaoH2FRSFWnDTd
Z9VziktR0MSIXQiutFXSZlt+TmcR7D9uC34gO4dTqPJMLUzYg+JtZpoqugk9PJRmUytGFqdeYRQG
yH2kxb4a0Fk/qN0q+pfyHV068xAnMDSh9TWGzmsogQyQ0kZqB4mfyxwuCieOlymXlpwU5s0eT7xX
j9eDHwHGQDdARtmZtsekuZcgZUJBH6bL1rrHFYR0C8pwiSjp01mzRM1qUMoDVc+CfeueAF1JvtwA
8TBqIiqPNENRmyxIWuM83DSviNSwS7Y819rxJePVQSK4AmFiTj+ZGUfRTm9HSz/71V7g5K9xOU6X
vBn0+C+2wGXsBlDVD0aD1qeFV6YduSGwoHy+I4rbjsbCn51cRjLsCaE9eTN0P4pTNPKVr1dzknKF
2X8uI/4TZEfF61cPw1uu2FigUnJy1zl109oKNoOHyr2+aSc+AVDt6ZtAcrEXYcF8gXwyJRGoJGrt
H568by1m4nqDlenV0cNAwA29yH5OuUcLHhQjWhLLNkKoDXIh5/uRWL/gtg8ieGZxEPpb7uZ2C8vD
8fUkFrHUWx8nIk8LGEb86+tR7jW7xeD1nAIiX+8K1zpFFlAsDcvzqbkRwwWbvFbIpBQseoN5k2fu
NOA/L26QYOatV0IvP29sjj2mOIe1TGNewteNcvjsVfTv1+h3XgcJUdLAYUM9T6WJBmBDXrMK1i8O
H0nq5KUVvD34Yk6MnujEg1WWDam2RPpBToUiyNT2P6hFy8um4w08S9qTUVwUJnTsJAGmYU4N5gFL
GbSZ5PzSK3kGsWsfdbTvNe7oMEVf6VrWVbuAxyfL54DA6BY6GKRj85Cszv1fs3ABQLDP9qf3jom9
inoNciuPj/nml4dNOPbnOXxrZ3X99Qu38se17nekP+eQ9fZxy+n6vL52Ai9K1kixrYvTjgW9CIdi
RBqd2b9Hh/Pd+0x2KpC/H32McjYOxvjJEp10UxEW1INhUU6qId6TPL/0BZ14DMI4zcX1fmLaPtLy
lNGjUOzHIhJme1y1mrFHjNTiwc0hEi8o8OXHtOHf3niude4Lpci7EA4XBB4NuS8mnpiV2vwOQhMx
pyrrPY/uy/SCyXhTv0Zx5CuXzkuL87WSE5ppm+pTwMb7XY0RVM0RksodYtEDlljIB1oZ6uedctU4
gvc/WvKln1cIjcNCYdkqJ4dKBTTlwt6NnOPwVa+pxWn9/EnGMgEAcGzTk/lAFo+Hace3iCkcJLhD
e0x9Y0FsAAU+brlbAyeKx8sb6+soieKSbSJ/p8S7VJAaFlUcXXn5FGs6/yThitcQRxGEyWfFmNt1
ddo+iJRr1s+u+uTA4pn7m2g60dmFAcVxmAIxShHbztZj3MxGqeAq2Wpld2OFfunYQNfZjxgKJKbF
2d4GSClgEcR3f5yU9Db5OQaTpOlv6ZKx+cYKBdyjR82AF/dJ9CAcyqN8ww3Dfjl453bT1dvRdRdA
78aH+RpgJ8IQbTPnixcDS+S8HgHRZ2XEiJEZgVTtbI9pTJE0wBEo5y4QE9WnHO/CWbsl6PS4h6mN
v1w/oHlYJswB7FVLyuE9pVzK3ZCbTwpcd3VBMsJPF2+gHB1mYHYXnQVkT1i3y5pPseurXWItwdvn
IsNUMSPoE1dMwzaSCjGSUSVIR+pyTZ4De8gj/LQ3Sw/Pw+VxRjCrtl80Eq6lt9EM7ScXWAHIabDg
aB4fd9vAYe2yw2S1gZGLNqGKWkbDg+1zPDrzHx3KJ6X0xA2Kio2eN/hiXyhoYSsNUtrWMKkdQZTh
ZzfiD33v57u8L4x2RxrExgGN5kKAVmAtgSp5pjMnICOL3ECQT5oP7dCnK4wCo1NQVAFI/Dgl8rlZ
bloCaQX4mWvmi3+En1n+Bj3NOizaolfvhGV+Y7y9ASzUmtOQy9lRp7qnw/8stWia9DdNimcuvzsJ
X80kKodGb8wjCtvEA0JuivpGb2g8d85KDy9sCpXdheCoghRnXBLZhu7Iy3Tn3AWnMmQjHBbTAqyB
2Cg7kjCZRsJCEz7onrbsBgx9cw/LtTJ/DunpCJ328PGvJrWseiBR7STC4DISLYiJLUJVPDSvqJrU
EywC0eh6xCotnFti0sdzc7ZThYWhQ82wxFDU/1eBChpw5DF6h78+QnkMXkC/4wxXDsHPsmL0qij3
iVYG3c/FwD+pMbeltwftwuDVTfJzIwX/E//fXjU3QUc/8JnuwlPk23jg0QJGzfuaj/Ut/f7fCUvv
m7Ec/vr2AfhzGpwJI+DJdH46cSHqg5Vy4tekcF1Pzyyp+MM4258oO20dpoine8ZzX50gyNVnQkkL
JYNm/sLgOrg7LsJqrZSfhtwpO7XaPCLVY9G0jQvE1zPEaKZOy5UHtWiiA35IBZQhv4o97m3NE6lZ
X5FxSmmy1tYPI7ZuQbQiQ3FTiGhnINrcwU0X47386zBqSrjeWB+G7Qb/Ai5JCvEFHXr+NSGs5x/z
Yj/rNuzFrAITLZMvZ9XcEEIafQupJDXwCqqqzshXYIopi6l4jtwUoUPVvBfaw5MKofvsy7Hpcfn4
yi5fErsdRcbUGe3Slnzb0W9oTrwsSXA/sbTn+0lN2GoLaRtcnS8s4NVozCv/09GUnQxx7KnmJOTM
5F4sKs+DdO84gnnGgE0s/WjXGp/Ma28s2eoEYOKBIQTYHh070A9JjEY+eO9tHa5UI2tfxGmoNIuI
S2SD+bgKITFqWLh1HSIb0wIxbIoKq0nw263IwA8RlipJmqF9e7pu4ucxbwzWu4hEjzndrohlbWTV
v2rJy8S74FAt8+4G8Fk+5hBEeVA3O9nuS3MPHEKbkH/o/B4/SAi9NuW8aZLuhSvrZ95NSz1aIzbq
5H9loLKjxHfX+W5EEdosw6R4UInn2H0Gay1VvUaJTiWYrRZi5OxcpyWOOnJ/gqPnG6f2/d63H2W8
mgHyM8T696fJgD8/jFKTELKWTyKwlGvJVRF4YawH2JYG163I3Qn4sTVQlpi3C5ngBc85AUFlIumt
RUtsA2j7HrB2elh/3oKogbngCQnRqE4utE9DmvdX1QIi8Q9r/sed5BZgNx00yw8hCH5M+DsUYhok
ZrbTetEUm6vRs454QHfSNn2xG7bbmrqCgFnASUtTDGCKXTznVQFr7pjmIaYxAPCLpwXYC5xINSyA
sB4eLHWX6b06Iixsqk98Nsa4SBj82RgrBoU3698amogSpBdWc9MmZBJ5uH83esuQKgJ9UpmiPPqg
cgqBPSmeQnDO+MUDdWuFMh3CAo/WkOy3og8aCAozUNE6QUU0ZkW59qn5jQ4YOaIOqm4QgMio6+Mk
84zF/FzGUONZZKrK0P2r6drgipvaDlsxHutfgrGPGrJzaJ2eFqEKpWHOXDThdFsOtd5DhtN/tP+/
3t+ELb+2r3RkblRpwzR4iWPdo7e8BwKlyNNYBjHxUYt/WCgeVv+3X8q5arzTruigGTW+3ydezB4N
kyCM6S3bQSO4AogWzBMKaZJaMNwP6Gi03BxIHR6iOWXxrheCs6a2rd1P5I3dzXX5wlb6F3qhzPpc
Vlssw+652xEaMgT/4Fy+BAQU3OTBvzH5xqezrNXY9KUHp6Oe+VHj/NsFyjXxvuuE3zylIHohDc05
ruzSRUYZ6di9MNjAwSBiKsW2GqOOl+8V4VkkgJSaDjLCnfy+0hIolAP0c8nRnPS2LleWfEsw+B4t
ySO/dv+mSlbDeIeaxVoS4ZYoieFqgCEowxWh8c6wsINdT4wtVqRcVUiUbxVGilvsILgL2NEdPLFu
n9/IZv6dP2XY25nKuA/2a81Mzd51KR25/EsDdawnTyeJ3SaeDmhNwHj89Fo6x5/IVJ/CHyULkwJd
TUzyQLanfQ4ZZJhelQhlHT/2+zQzroOm/NIMedF4lIidOCFroNDUWmV4FLSpUQ2H5YgNG3BZX0Yz
Wdbr0nf6P5j0trDzZ3a/g3eegDCb+V/fg8i1agyVC5f+zZ6AFGaqlvRVOXHCk/zB+uL+Shju15m5
LT/63izW3ToXtaVIAVrHYdQ2VT4YP3hPMvHPzdWLmQcsuTiB1Tcreuj1pWSzK+BwVqzZpBDWWJZP
85e2rn88sOtjAG9WIrMT20cLpNLaMOd6FD8w7G4kUkyFsYzlxnYSBdwfMvlSLr5m67XKWXb7kbMO
iyfcxtiym/z9i+9PBP+qiD17j1+nGzNSryAv8+aNd8a9e6IDuEdghasv/XKg9sx6qdggo9+Qsh+w
Yz6vHvgwGqJ3u8uZk+699LhS/piEnWNI+/Lq5PgVMoslT3q/VPDau5rtbD0cyNhV7onV8orD1omx
p0+p1Tn3S21OOmIxMBFj19VlteuyiQ5QZ8Wb0LieU79vRJ9NwWnVQLslJBrdFUzR+skU1XkYOVis
dfwRxQctuRu0p4wu2OCMjCFt/Xrn3805F3cik7n2rJKbabejPbcr6aZbcQAC9V/uFov6arROyJCX
unOh7EU80Czgv85j92yZLYeuBR2TrU6SZYl/xfWWD4koM0ULayoyNbEkrIbiTbqeb95BcZ2f8052
OL54TDD4+jFnDT/mCCvihfAc5Y5Wsj0pMevYQ3QGsw6OHTvJe6VYD7clvc9tgsFF63bYT7oUK2GC
Gm9ZimYSW68Bow+0k8vR1b6dBy3u0w19jW/kvdCjvQumfOq0InJcLfjQMcqwowz2ia1UjSQAH1pi
7lCg6zSKKbkWhNUpFhU0AX2sdynT2G91M53tZnNj486lznJiCfbQt03iJGMqpRaRmgCJ1HTti6pC
TYt3aFjAXqU+H0ZygiKFrzrUskBsh89EppydhEEtn6Yp493sCdGQQQFoH986Gb2XOKGf7kkXUjrn
j95lR6m+jY1TdcqVgxu2wbTLQ18wMlIVdH5U+rTZlQd+KMyHdMTQjuMFzpdFz6XB329MryASOMM1
5wKB0GgruphSdOR+oKORHgRVKS66TwaWw37fEI6IrdBMNOJcH0dirmBpmZET/KUKFhjemR3iRck7
NncDGuflAPFFEerfpuS5HNkyeYtXKB538OnXe8Qyd3F/4ZMdRuBGtfC5CTV1S4ZHmIa/+oa+LfNS
8LB9PT8k4AxECK18l9r0qNpO1XZy199A4cndt/ZsoeNun6rprXb/C64EQSKF1pbgfZ5dTl19Q6Jy
RN6FE6pf9Pc1lBrUw2Kpl/rnmB7O5VWwIK9mvI/JQNTGNxlx/gZOw2YRI1zdX+j+lug+SCCPmUxP
VCXCaqwnAYgJo/r2dr7Ionn2n4uT9RRJi9xQ5rRyVBkWkejbIIioXR450NqpzhpelV9LHKKw4eS/
Jk1yJ6iYoRH5KqMmqgxPyo9sNWEAYyD8mfEoBoj3EvjIE7ggRjGW3IuD2LGsLhL91kWAsA/KWxsN
rhLTqWsx6k74R/HJ6uSTmKPp8o6AAAM+jsvyRsCUhZEsRU6U+7uimS/Mr5Wz8Fz1s+l/YVtyAFPK
RYoSfnlr2/jW7cXQxujQC0AM3iVyVxjdkG1eHNbW4Yfpwgs9kPoektqtjmVPD4HdZaJG4F3/8Iqv
caTX+xiTzUCgcGBjQ15DZDERO144cyaH/ZHY0vfV6VHyNd4oTqQMzTtbSKWAQiCZWQgyhKh+EPZB
XOj3pqpD6lKlI4XP8nkFIo4JTHk+N/VvhXNMdHdcyWqBamqgiiW9x5WmfGknoKko/0Otc54EoCV2
dg3Uws5bxAptGKPBtJQeeMDHF1U1tbugxXnCJFUk5ds1wDl0ln1zrNwy2AohubqiOn/b6dr0Z9T3
aiTNYpqeLVdOIZStcR46i68PCt/JqZuHBUqN0H4UgjOS42efA9FCymQT1ugeDwr8APxyQb8nvMWw
6pbqgTyQBZeQLkU/IajIt8i6pBIQsONM2BN7Z347hhV4sR8z2gaKND8yMfeNiNttVoH3HXdUDAbl
E9XhuebI4qLi1MZ4gO6etesghVPB8cb4hv91NJhyzsG7g26f9SPW07fOUpzxN6s0ONiQseYKWdaB
AUlNCDwIkRv1N5wpID2XznOoYLu7K1aki+6FNY8jawvYRFGVuwr76kFfBRmZnTMK7bf+SwDdNvXm
PKe9MBqYCgKsckStzfSzU2jIRFdG72K5Txfv192P2zaGQWOXkxtoous2G0eZesws4xk5hLlLAdUV
lQeppIdfdMkvnB58ouizf0cB4UW25D1uCsLIIX75nUXgR6Dk6SAmVmJMmHSbfkCEDd8OIw6qr8fN
EhhreJaNyLhyvuFbBVqvqk9FpdbA/QHW+1KoBrLbBX0JdJ6/liwqNPTkKwHoGMtKi/LW1iiLWKuk
CBBQJs1avBLrh08tf21umOSrc0KOF1yq2CObtXaQjX4KFDOrB4xOH92Liev/Bfy/uVcNkNM98i1y
3ZbqeRhsOidmBuXwuX9GXmuny7xg0Vb0kryWRx9A5XewYKfVfjfpBTueX/51qb6xeEO3y3N7YR2M
b/eVUmlDfy2xaQNCTZcGPmFc4CxPSyKHpX3T+plrYhckQCfUcn1mZU7zkkCFdOIebiEQrkiJTrO3
SnU+in1eSI73V5SmxFO3BANPL5j+vl3n1tLz+0u5Gbbcmq7Okqz8P102GNW0rZt/L/SH10PHYPTq
GyJUB/cHEi3eSY6GUbcMgUiFvjJ5uxQJI/+64WD5oSEKpeqrS7mZkQFQzZdTmgyQPh1r+dL2nwZ7
4pYoJz8sSSPBnduTmfiMdliYZkYpCYgkQYpEXYaJfE3BrUMfl4QqcYeidgTPoFZvqICZyMDaO3Al
5B/suhcseId0M2MWy5pFI9/+rXR765/RL0DLg8OIv6YYpyiXCInTKiJLI4qTaEkZ32mqFJz/sSSN
h8CS5Pb8+t0IGMjUoJFTxBZkIbH8zed2qMLTmCzOddHinl/oikO9hXCIgCE0Rf0GaSOlieKJQVG1
0IcjamZG12GtpEl33X/3GuES2qhIgDzVRICbydWGwfxOr8S0WlRy7Co3EHSz7uGU+yQ+YZx3phht
pHL5qo7l6vCLeZvrgSXuUJDnq1VpspgngpxOj6OUldjL6gScJUrYlLVI1TFeaJk5NVfOyQSSq5aG
QtzpjHFExXPo1mfILTHa/G4eGO0s7biTuvRxRzHRG8ngTNKdwJ72Cuv8QP656bS1EuLFTomiUqkP
4HU2V6ZP6xi2usisroaTmG8Bf09VJY2V1PuD6HAK0CEeseaKkjZXb6fbge9dNHC/igk5qhNcuTHM
obBd5pVJ+6kG3h1XgWGhF2/w8WeL1J3g2yD+U2LU2a542GW57dj8FCJyY/tKlIAXRm8bYh/5aLjA
zcTysmRLkop88Hbh9kNi3iBJKA/YdU93BCbGHI5ksT4FAdTn7dM5u3yRdgVPTpDmr1wmK9gMqLsQ
YZK2hhrKph/OXlwTAq2CnmSRlp1rWssO6Q6GJTJ2oVNJkWTm+CQLSaaxdxHicz8zKu5a+/frZqTR
0otD5X4CTlQNojQ4lzB+AWo8cBuv7V8fWdxMgbXA+AToNiCXVL/l+1TDGuqsVzaWiCgnOlKC+/us
BWrHvROS08kw8H40ZDDzZt8dxtio4qUGfB3+Mad61JK50XqE9JYyJxH79HODcrL0FwDhbgmAR455
r1TPQ64E8dCtCnGFHaH5VGIknKusViG2bQd+fJVIcLMer1GRKsRTDlNSpgi7zpBE3nnIQJZazPvQ
l8L42aJJyEp9tAqW6JHQJyt4PCJHLoVUWhituqvk7PzH6spO4f370FZE/WRMtPsUF/rle6UgwL5I
x/G3TEmqtGHdVMuptYY3fBA/7GnYA4FEZDhWPHxWtjWWZsnbVhbp2L2qxMJ3dtbz7nM0PvGAx9an
hWw8DrpFjOl6YVKLRT1crxwIAP5clpZnesNOCLZW6TCoTNpzfVzOsajy8apQceR9kZK0RzgiUf7k
/eyYtj2oixbBNkZPzXgzcynBdIVJzaC4hLxNXams1FOUn9hNqCEujP7ROwIatZzhp3NKMbObcEur
Td9CPi+7LbeiW6lRRf4iO17G06w84LEoWyppGDqjzr4y32jCjhf49pYM7vH3NvSxK1YnYbITkptn
MjVvHjl+KiyWvUA55xgFF0glwXvfeuTtXJCemz8Ut0o/70SJpeblHtGzFEWHvexlpCrZsi4fUBZt
QDROzccLMRjsKlrzGSaN2j2wJtxQN5j8OPyHFW3FglCq2pUErdF2mxl1Yk56agJlyOEesXmqkvzF
4qgMCTpwiC+x1w4sWyYci1A3npMmeDKmYgN2gGhpOFUbwSy8+QdTQoiuU/liFSTORL1R5wmVUxkt
qRiIWrGKuCbeM+1pl5VhAts7UBDbRZ4Zml2bcInPqiWJDbZBw2ful+8kCNDXsYeQk1l8urXc1Rju
hUFJsjmID6Xt3wzqdQrCwMIy9n0/2AOLczTKNcSVnQ3J+57B2UKFPQpKnb2RwkXY4LXNFrD52Um1
vdSUlF416p19VI1WAYMpqv6NaCuyvy05OZDcR44RbG9MPcQ8dkFtYveh5ATHjg0rIlhwHE2ipAH7
GHEDWo5bO7GXHRVRVHLnwZdwods31L+duJGVNhfsYuxAWh30PMt5HiM/HNGg1eZLH81iabZ3fD2I
E2boz7TzSLpJD1Zpeonp6WaKeEdVEFp/xwGw+bnQdV8Wb/zyLYx6Bb85BaxiZePJsTV40DtDkSRE
qqo3bk6QBenTCRpNqVtYDWzoTINFw0SkyZOpFGp34QU9GcOaFMBYTV9U3RYgrLzm9I1lq7/IpffB
KLMSy3SCoqb5uMJ2AS+fK9ZY7jrbLrJrTTV7YWnTJSKox0i/jI4ryUJ+OGx69YD4Jgig0nBOP265
aeoBkQM6wQsbgZfpXTvsIB/qB2JSUwTJVkpWoNomUsoulT4jHrcZGOVt+4P35u4H9tF/M+QAJQjh
I5wRcD0/k2z51tq1YO3OXsyPM5wdq4vBgQYUCs9Tml0Lfk5AFHuZv754QQw4cOEe0tUrhRZ31D6u
sEgv0xLNOEx8GJeT7tJXcbby3QdhpDHr3wSdvTzHs7hJcBTH9xJ4yattqkHJPcma3JmfrDnQ3JzH
P6y6HYezXhJiXLHx1OyprGL004tPpSNbY64xWG4DSMoX9nVN+xC/KPQpWKdQjj7uEr5DDG/JPJnY
ijcfU57oUJC8xXGMsf+sYE2LQ+pKeAaQm++aua+clwmTvR1jYxJfN6JX3xkDCIfz9hfH8u2bgy/G
ISEfKdpxO95fddZUwEHgTMTUSnrRFQO6f2FDDym0KR38f+vPxD8WBSq5FT0l90Evxb10nmjtHfkf
jdF6vd2MAZXtZT+0FrSji1jEsCHp4Fh2dASzshEKJaGns4QT4kHRvYTSc0dVct5U1Okhcrv0/Y3a
mAM0NPBsZyut8y5nJ0PIHYUr5b8Jn/3lxc1/0Isa5dFmFO8bSIpD8a2RUwHpnTTpe3a6ShKewGNR
ufw+h1MsCSIq84dhloEfumLHZtCf5VaIhi7p7eJnZu29NFnRYViNN/D1wAdIeU3aiyS3O531DH/O
a7L2uqU9pcgoCtUiJIV9g8W2Dc+qUx88rUZVgKNOyNK0+IbqNuvzNtJiZCN93nCa3eLeR+FccPEm
HSYWJHyHAVohu/yzlubuYm+RGaqvpeS1Ob2HFpbODqMa+cgmto9DFd7TJLEnS2WuJHoX9Fk/FsdP
FiOMWx6lC3j4QC+/ExDI+2cPvNooT4ztwZESyATT6JTykPz+oqyOv0tChEmv7iv1kEOGVOfszi5a
eAvK/xp0IiD0GkcpQxpxr20pjHFJOHv1bb8PvwIB5SapBnFuvLFfauP+y1sMBg5WbMt3InaFH2+n
9T0b4oofVcEq3yMnlmRs/hAnCK51K/FJRtBA66BgRt6ph1WlnRokR7Odpyd5Fq4CZqsHxwhRqcoI
aLcQ2R+vLZePfeNfK3etOnQHgKwzauA3UhUwHyUG02ggrWhnryaNmG7iGT9WmmCoKTQnsCnEr8gk
yKfZu1S8fGcGuSLA68nnHLrigt1+WfE7/2UP1lXFX/d7wiIEmKTKgDi2Wm3G088rg/1DFZIys//V
EycljupgvV5UyDYxp0xdjQOpdfFYUuhqdYLUsNsM69y4UEvmrQF6xF7VzfXoOTZicjTCMhLeRP+U
4GZnf7oKFF34LedsW23Q6hr1SZeSlM0yZt6WcxaT85/aSkYnkz0c2OoakZmG0usUET6srM3MUkYC
ZH8D3uwrAPSpV44jEvxu8CtNw16ysm8Rml8r1PxPp4gwAQomTsG1ac1b2D4yr/4VGnEYXtZjuOPp
PAvyTbQ8KXLWh4muU6sgzU512RgAagvBNUfogP9waVqwTs7vMsdY5Ua2tp5BFwxV4RKdhfhwjAG/
iASq4VeJs9BOf0Mch1g7BgB2CEk6E9FskY8NSXxEdN0+JKAUoRPvG1Mk0RcbPYgi1uIUy3M2uyvN
7l3dyNwgyI8gztrvsNNkNxuKAr1f2EHBxJBfv70OLQQNbo47bSK8KrKDxt+Ah4mEX3VWMY+1hT/5
U0MFRkwRMUvIrjJQsVu6NzfIBzxMx5osI5sRdKOZi9og0UQxPfb+Q4VBc1JrUJTUyZmt/2ikcJBR
j9iBah2blB1CXw5ZsmraPmKBxgziK5cqODGzXsvZT0+3gPI2oSwdxA9FKfu+I87cbKgFyc4pLXt8
sOo/OBG5b6sK+Af2vJR8BjPXkeTnrM3hPhsP2WmdM6StKqmvHnRYREcL3DDpWDu3MhzrrpFq3HhX
vkw698Sp1Hu8Rp8b5INJBtRsen6FN4/u74PLNaAlzgJm50uP36HYQGPkpbRRZDQXFqMb6ZJBlsWM
iIO0oFY3zGK/wUbEgcm3k/aKeyNAXeITnGXTm13t+7OXx44QdJWIlXc4WGTdWr8Z5hhrpnFDaqAg
TtorIrDnrTaV4Jhfauhr037SSNTe/9IXAaGCy2aEifoPKjvemQCVV4SxX3EUb2VDRwqgYjdeYNsw
cETleNj1xAqvCRdIuhX+uSEPFIEJWz85qkTJXvxCLnawE7tW+HZv2auF5qRlh+XaA42PSg53J7PL
FXcEetwnnS+0bSAgHQXAJ21IiUR4XW3Z7Qb56rzFcaDUNHZ5FGMD72a+0PDkRp6ngTwOjvr0FfxX
qsFt95L3mq5JYNjVFO9evaEDr/I6qhdxfTm+qMG/XYgr7sMEI2YYQla3U0klXMrGgr2jiAoPGHXk
dnvYfCnZfY3rhD3z/iX1p+ZFXlzJYxznlAPbi4m2P0yY20xhxCcMXhv6yiyXWVnsWrJFaVsR4q6f
UCN9+NZ2dbNZFQ8wyetOEcY44D76QPMzpCIgHpBbIcDcXlSZQK+SbqE8gy6xuE1CSP1E9SHqklOj
LFFHFoVZu+/3lj93McCpd4f6h7nDmJ+WM0Pq8DeqMoiZjVv/sGt3yTFuzCzxbOqLWa4+KJVltdti
0qcu8Ylrq3Z0Ct7XXdru9S4pz1raXby6WwGwlsS4nIwEidr7h57M5ZkW8GzZWUErOpeqzj7NpFkk
OSAr4xdQombSlBsKEmz7X9ohroCbay6LRGPacjVSOaMvbx/mRK2iRyc/9TCP8gmjNCZTgmVcCjK5
zmTFTaG3o1V9jZXqFzgNo1ivFbh3bKzDOcTpZXyaQBQVOOxg86bGLxFiEBRwmX8VEecy77dGTwj1
D6H1KP2M+H8RCRZ/wLfYb1R11DfxEtKafuwV/dDJyepL3yMqr/pzbDfmQbx2vdOgqkosUZnEfCxF
hhE6YGD1zbumj0lU3fNzdIgu/UuIeklppOZTvePM7o1Y7et4VrvpPW6OrLJ3qaQ52B2PNDPt6MDa
jRY7GuyM08yIjsxaljV4gl5MGoAa7Xk4bGnXSpi+nk9NjiCWDhRzQ3THdSGjcMCvjlSuHW+gePQf
kJbizUEwNRjL45lCppVbO27m9Nili1H4sE7aExlD63fL/uiSVyRabVeFJfFV9QTmoB51Q7okmCKn
VzJOJ4JUHXoX39et4ZQUiwCvh02/Mjh+CG7ImnLyikOIa0wPa+q4FZQICdmkLP3FoWfhysgNt2/i
eoEK/A1HpVuvGnrWV5oyYqj4Gej2n/MuIlu4rdADmEeOqDY9SpEaCx3nOsqQf5PYDT6g6Tb0HE33
GwMR1Mea0mmeGcMTZZ0WliXmOQq9G6pPsylFmvO8oKbjvla7s8lCWItLuT3HJpKldXJf7GhWoWZ6
wSMmXDQMYsONyhsUorR93yvezcmoG+iIYkpiBbKUKqDXZ1JuFVnvIZ037oKRrJY6oXPKCbEZm8K9
Ui9AxG3byhxnmrcFRtnYA1yk6VW5w+TabdNpozhSBlZ2n+6jGUTDU4xIg5SdwWvcisDVLBPFfD77
cIsUjJygsG6oTggiahA4Ewu+NEzbAKggPeCx0mgivv+U2Rcqu6Pb2QxfzW29+mGxR+VELGXl+nkW
LGKwPri54Klp7dRNDkAB+AcMrI9B86DJFIhpUe/sbK7j005ymmMK4L1mTgw0suU2/GCj2FZaSyeZ
NyUry1hOhFHgmgAGIhcvLFx00FfMljDaLdN/+5pj/NqlUbhoVrgnujuzWsi8SDTSWJrmlnXNDGRX
t0fVBWUypYzs87bVfCbwFN+ri87ZnwCkHDtD/G/IJA1Y5HB/3AdPMUy0mCy2xiuxjjwdGXdwWRf7
dL2Yc6iNGN0TEgPH+OrIFrvwaX7s9mLZAKPvOh6EFk9hzrr7l3H/NuD9tT9lAzHRBHiDPfQeerBM
ULSbsLNY/5rAWTfhYVan/MgdTW3uyXczWqD7XFtMuNpUhSv7t5wMY45bXx0as/FQWdjNhW7UVoo1
fiKowUniwET62gYwR4tMnMTURVdQhlBd8cgLeOd8+2p15hf3i8rTnXsncNf4uiHpOxJzmGGj8two
+jbgVE740R0GD8Dq75jFqyUV/AMfzkTEJvnRZCNpZcM0p6TFnrrFRgO4SOAPsGnRvaf08yso/DOc
56M2luJE7q/KDd6C371y9TFgskEFPIF3o4PEAfyKhoA6xnI9VVYvb0w8FKdrxt1LtWxiOTBbczPn
vyB/SiL+DO8RH6fQoGMK05qsWDwJEjK2p3WD/MeGKsCPL3XfCqRdJDvInxVEtTZMaUe20H4q9vK/
fQsSYUCbURakPd1y3lONOnr8enq3VNWy91ut864vi9v4SDRaolbp+fTkOkJo8Gqsr/en7ks0YDYn
s7qU1jLRiPRkscjN86ZDioTD2sKmga8PUY8yQjL6Elo8666wzGMo6mxmPwiGd7dIhiZ4wI2o0OKV
auhUBhtzsmruYa6zBIIborsbr7DuBR/k1f3KR6ge4ijioxjeHydp8ZT6lwQPqM8paA0GVQFp9JP8
wQsPsFZR2Oz7UPbLbdx1jDNNVOoBfBNtMry9Ke8YY9cwyo2Sp0txNryZ/eIGtJyBadcb77GDTknu
lxcye1vZfT7Z5eFS3/w4zitnwECimxtD6YTKMUcWk5lo8N/53GFGyrC8Am22ssSYh6x/YfLrIBBO
tb+XdzGhLlgODSYJzf0snO7yoaThAsopTOG0ZKvCyyPPSDD/29YNE8kAwdtRpLmZPU58aY5PUqun
WJsehoCo5n9BR2fr5I8FDiZMaFz3uqsNUpuqH1ojo7yjUd3B3PKSt11pPuQcQ9dON1PI7lzCgobz
CvvoMlDr9S9nfJpE3U+rSL3JNi216ldiJFtUt6PN14XcAJT3fnb8qJx/HH9/0aCsqOVYnubQifp5
Ikles+uaSF5yms8Yc6UBTzIA+TFWqVWV+QB1bpHwl8jv7EJKeJgHCSYDDsEV3VSLYL9YOECh+oCd
7X4pFa7vXj9V80B5PVO6PEjAv25rUiLl25nuh7Nd2a0Bntf9yFtIKKTmA3s6XwzeOtyp5ZA+4ukJ
y124aEAEMJhWRnWhpPMD0npAovTzE0Pk/oGsDqa9V5rHbh0tnOMjD7n5cQJkB35YTlo4ewvZWU76
VRK3cPxugYipmqsF5jeABUfK0HLTHPVN08yl4SMa59P9LNB9t76JIV56l+zmE+UE7UgevPB0eKpg
hHDbaVk3Q8O7ORaKkw2Yo33IThs0g6YfHUstaqmTspdlAbzCWhAyWExUh65pSSND9++mSiN6I1yL
L9qFpgkPOvVKBXwdbt/LHDFPeCGG4XTMUjCkYNEbsHtxfInn35fTUQ2VbozlXN43Y/V+H60HwAYt
ut4OfjiAcAkEwSwJ0WUr/T+SX6mFQa0LZfh+WwD/bQHaQYAR+Hgo0EmraGEp9DxMwjRdJIGpS5Sq
sOdI9vOawAuo3W5Hzd5mZ7AXWYMO1voVACQeIsc/eVjF2Qsvfp4nMXbZuJ4ItVQ01Ico3Xx/iBdG
EJbZVHLDlPBFwQHVd6B7baDUwfQcIj1btGwsc+ECq6QLpQGcYa1/NCyD2dMZ03NNKTxsavfuuxoj
tQgsPI0ACJnvnxQ/tDZHIFNbwF5w9iwmtr6L8HPv/KUVAuJMhyi/wM224rs+OHTXU46R8lv/NP8F
bMy6P+3ZtO7N9kkTTHstvAYBPdtf0M4kmz3jEAvk4Y08koX/O5yTTam4ezIcRc+RC+H0G3eFFTi3
HRqBii9ztXzj2F7o5jtPbzxhGLyLp8AQ2aumF56WGH8kJLXgxGau7nls3zgpYmcyzR3oV7AVExHn
SGZHl8kbbN4jqGCyl0Yb+4ZSyOIY580t+f0B3OLBZkF/zv/SIuAxP65EqyYfjNCcZvVRBTGKSYRK
mXfm8Dz/aCdJfQb92YaNRsW2FD9TMWI0rAUFOnaYjReD0fQDIJtvWJIKCxRkJ6U+xvN/MrUyGdG/
McbsuZoBBIaWRGiUaHSA56NKepvGY5ZX6ioK2qQrpgloNL6BBdhVoSBr8mXjQiVdNpCVUizqy/a3
2wBWxVTIbE+Dryf0zF9V+pjDCShuXKZTtsYq7jfDNpQg0BD02mKKC3MTiZYxq/M26L7nMG4i8XDq
mAqv7hAlh8ZWPeSRKPYR+6Z+MzA+Amiji+/roqPpsi1zb7fU3X0i4jZTErKgHGsWAB1QRt7sy3PE
Kzmlp+ansOA517DTK4ZKirKzEUdPm6y3HfgMZS4WbGirqOLnxgRSo6JaXj1DSma8I560shnbKcFW
6gyfL0eJzmDWd2SrDtLx/MYB+GW4Im7Cjg+MxNLYbGH24HCTiBZwr6wgfdFoaxRp+b+YL9xmGgVs
uB1K0wReC2U+bQ6D8VRRk+CSCypmSnXpkq/Zb5yL9WDBzl8uEKAiQSnCVyL0yGXLd1yXCwy/3+KW
h47TGU3VtFLANhSRM4LVkKjLTFExvTdBMA+/kgbG3nNzI4qbvzj2dsXXp8JBbsh1NiKeNr0CnvuR
UwRROpNlxvo1xDYGV1SRrfD9Ny92C0MAaoQCMx/JgevuGWYDUrO2F3sk7rJsD/7maVLzbIbeJ0Oo
Qg1G2c4DrBUnNPF4ULl0FNN8ryQhBbTiZRswBWwdX5TiATs/sJEjhceB8gHXRi4zNRIC/SBRi9b5
3izgMJt6xQ2Ri8YBqDKm2658Q0nUB7Y9biRbdROiM8nFahp4BdyBAjtH3LpTo5GRqPtclMyy1van
3YorLxOvdgF8dqO0xE8EnTKYZTk+OtCgsfmqgfWl6wK6XLrCwrGzN8CvgoEaZYjhSEr+93P79trw
M+xDJPCeVL+kWYQNA/jC6McZ30dSeF9u4N4ttn4DHPsyTBd7WlSui7AvLFYVqsUAlA73Y9iNeSvm
0JtIGAOz+WaxjKXn0ngFHRzX8M6CtdeMcfrFq/QHY5gnF0VnfdKsSpvb40eLXuzfXY6u7lyMvfUe
74VgXzQOzKpomiT/4Pa2zxtu4uOEI8u80NXKYfQFW1zfADhiYdqcZyxFPE6tIMCS4dU/aZ5Ab9DJ
9/Or/p8x4aQ2HQk264Di4KhlxARNAuqcqxW6+l53s65ThBYqdPlPeSBYPtQ91qNliW3t1P33/LHF
t4jhGIcu2pdU6tFeJ0cYDU8kW26LYfTtoDdhxY+6gxD7y5Bn7CU4mch56F6pxK+Gnco8QIN0D7F/
MUf4r27QdYER38Bat0kXhjbuHj77z8IX0WgjNCaDYJN3g3FGgU2KyF589XsvejWa30Jm8e1hSyWB
mgoOAAiuqKTD+I4wzwcYvEbp+MrXcU1jpk8whr2C1nZL71s21bNhyBFHogDjPoPUABrRY1EXdQSw
gQY68fGjdknNL0UPS/70ZZrtARcpQGr95v7e+PTx3pdkRUpNWpGSY45Da91KxnIsonUslXEOZXGb
vwjU3ZilhZ0iaSLExLUW7RuuNEUkbpIP2rlTpZgsufc+43hxNSTkykLh1vUUIvuusdBPIqqUP1F/
ITNCVLZ6bdCHwdM7sIN+1pZX2cY/x8O0UcWNgZyFeb7vh8ZmJy22Rmy6QPSdMeEk4FhJ3tiZE25K
ZOvzzGghCw1anOwL4aSo1j9j3nC/CSlmRl7Xtvm+DlcSX0QJn463W37Yln+NiIS08/lAWp1vli7j
DcuNdn9tpBow8sc6OkEhk6lGP5D+0dbjxONQEgMnmaB4c8Oqtj81DwwRyF55ax/bZFOJspfdu+OW
1Za70I5exszzSCN/hCsi6q2HrwwbqC3lmH9FMHTf9lOnacAPSdn7Dvw48celg2Kln5qO9K5lqedw
K2lwqEAiNZvia3DR78LcuCo9Q/pz7ZziXtvH+WOQdk4Z2k6gDbg5rGOZw7Df5Cc9PbJndSrGD1tl
7sGchVTh9LPK+Zy2rbTGQvQSv+TohebwhKxu14TI8qYL7iKF1Ivy9kI2e5drYzxKiqwcn7bsiQGh
Mz6WKVBB3h/oZu2K3QWtawQjOSDQAkoYS8mdIdoX0j6+1LYxoB4VOO5CiD/Ggy7PmBCxlZGxTklF
d7nF7oDISZS3u/pQ4o8dNktvaR5aQ4gAFWNERT6OwO7bOjWMO0E6VWxlOPbSMyvkB7fUUOYacgnS
QOaUDMAk2fIz6VpGiyATxX64lBgByZrQkoGrgWZXuyuQF9dUvi1W8wuQqxIM54u4zS/jCUKtz1Sn
E5zFd29oJaLCQSTgoMUxGnM9vpRpAZdW3dYqq2R3xOt/uQJlR0igEDN87xn68HG7odDTHWrZctg0
JS0xsLXjF4IC9FFLJy3Oz+UWk8KZTHpWQdaZlUkWq+3Fm+OJoH85BdyEUzzEukoVDRuRZCSRlW9e
tAIinyxKG8pSbS0qkfae9yr1KXzDTvQrtqlD9qOzh9N14Ez5/W5dGDEXhbvJo/09zlv5bE14i2p1
kSnIFO8K5Dpu/IVRvLNpz0IIGA44T1eEUo/rOrgBHS+RONuFmGa73AymFBSQfrAORXHgp8yXiGk2
YC29IdQcYc90U5CVq8IPYMTrrZI3FCnKU4cfwMxjtB/zGNPs39lip6RUAMiEWuia9icmEL7lV+u1
IzG1vUCrVcFMFyKerDqeQlJXtKIomHfgLetZ54WVS0yi4kGiBAhOM1XZ8Snqx/ygTVBDd7RFl5rU
J3ezBK9MmyhtYJK0RQdrlFIACBp3OFEEDv0ovztX8lZ5bxQGqOwalar74GiLfBycvtvVgUIko6LC
ktbCznOjd35SbFAB7McIADUQ2Y2vS6RMFTgOQyx7kkxIRubfgDv9TdPcFcKYQTUQwCf9NCrJPWEM
/3TCev4AiCAAMbXn37uuz8yr814d+y+0JTDi0Nz1E6Hw4NWVMh2iDTN90M+qSxhCy9KMaC8LnMsB
y6wJfD8x1RWyD2cYyETZB1j/MNLKageTQnuGT9ff/M438aEA23HrqMfh0IIgtHtT/wxNOayW6deA
bQBwS4B9x2xTRvma9LCwAsjBUEEPavR7qb8dzybiUk6pzxciaxc2TTqcInJe5cmLmOYHlYoNe94y
3hxJCDzhZi4gZwC1/5FsO5F4cGjUvWtGNbSDL7uL9fDHg4lHosi1tA1W0Yibns/DTVZ1cUBXEOvi
r/ehn4nfRHru5JdeC6jqnhT53jhpDXWASluhNSFoPRFD8ectYwwHuYnyE1xHdAgRACzT8uH2JNxY
6CmOj7QszY9x/qwtwfzXSt7KrByB5jEZw/ci2GrPPB3aXqJ5Zx7tCs2YDfSE5BfpB+wJDRE/mbaG
OqU8frtZZ9u5kYvbR1wuc3V0/tudfih+NB2Ao6ap6EKAcRFdeXjFZPKpax4Dh9IATkbUG7Qw9N81
OwPLcccQ+a8tsTiyHCDpojXWLs/FcWXyEyAt5C/JAAALDcrQ/38hJMKKtoa9LfJJLAxzqSlZdMdC
knqU8WjsSJ57rwtxQHTLG4WFNFQ3W/J+7J3ElpGoW3KzmqYIVvNfJMBKlJcmOVyduysM89e8ys8N
IFJ3HNOVCgTYJiCNUOG1C6klNaVwK1cg+ybZ62v7/U4Dp38cD8spaKq4NkWvia2ZFq54Ssze/zdK
IDrRUr79qBf6J/AQMpAs3fpP06PhBZuJMjj8dCYBR9CXoo/5rwSeJ0gaWo2dC4aZE5jPRXIsKLo5
Nd4cpq6BEPf7mXvgyXSZXq/Zb0l8iCLIJ8m77FC2m40VDropSvf11ls5vMredyrMVGTW9NpBv8Zr
wtKCoIAW91TApLbAFX5oJvs3I9GEvC2VsVAODnnH10hiDp6JcU8LZF2/FkgO0TPzSeHHaOcVWXsN
b+3tzzuJowPrZ5XpDYvq9PB3GpJtls9TsO6xk/VhZkEM09Cix4yDx3vwNAX2i6ZUA+w8ZZ5dYooo
PnNoq51j/pEsTu7AlfYseIpwAd16eDDN1IZJwLymYea8ioZr4ROGkBM8kLjiqddTRCGzPEUVUTHC
2XeiYEDwpBRoTa3AqXqwNCH6mMuNuU9xmrNYe85fpx6JN+eUgp+4Rpk0nlPMkmfkzwb2ulxITLjv
lmt/NF9OxtQtIkvafK/jlPem8n54wP4wX/IvnjV3Hw+IUfvSY2k0Fdi/XCdnpPPDvcSjl4Fofi5K
pkjCIbp5HB/eVWmize93mVgxCDUhrFPdITFV7hrvs6dMEUfUNGuCJHBntW24nMqR8mM6O7aTVWRg
iiY2LFors8/sDVzugjzYowAcbu3vKcHXUoBMN81hnQM3vvUJFNCwrIl/6UCzHKHoIL5UOtyA6xU/
tM4xv0636bk/esUKxfBtLitGjq65R7Gajl/XBoUIoi5HRB0/SgWP1dC1RVrNOlBthPObBHlXwm+D
ve215BKZqMJoWiOBR8QYK2YIIILL8Gf+2c9STxw/KW36trvut1nzEZgy5s9eKKGhUG3O1Q3PTU86
mZ0s175udoeQqw8Us38SQ/QTsJzDWZzz0MVJWL9kp2o3lki9TE+cLYYAEz4XFeOlkkSF5ZaGBRXN
KFqjHs0oNW/tNSdsntPI6Gt8F+btaIk9iABa1DZS+9OZ4U53ReJTcdtShL68tWsMYrm3is8M+iXT
RzDqYsr2b8FqOe5L2q12O4Jv0NNDCMbDkN2ZX1xj8Uh4WhOKlXdy5I6tB6KoAxJcSuzcy90chSiN
bSgZp9RxzALEVBOq1S8RH8Lhwj9FVYzqbi/YOgELsGh9Jz3YUvmqV3ezd2tBpvXRg53+z0I7X3fY
kzOZ+DoF9ACSekasNw/OmLj+YRT6d/XNlvOibgFBYalIKt2oziCP2E9FD2M3HOMzBKtbJ63skNwl
ZJOyRi1ahYVeaYRKUTdyEO67lt54T+rIqsn/ENEK1nBay3D3GCgGSVO6ZlVG7ec884OGFJNePBaV
H/yWCgAGsOUQQUXkR5IMZgmQvxoAz8bz4VDlaRKvrRr4BRKAvQbZQ+7ZiiUkxrN33CP4e6y7C23L
xqQOsTywBFT6YUUz3SSp9CIjUfzvDBa/K1VO233yl9Mibs7RlwSf9yrdTNls+kPF5dPkUcPQMrF6
EFr8A2XMR43NJK4V0lvD6L5uCq9M4zPf3fcF3L9TUdb2DtI474nRo4IXusQXhYeueNIG2APL/XNo
bJrqPp+qe2R9Au8zgmh78+tun1voupyhx4Gmf4oWHLS/q/qftmxSmxp24cQLmtA9HvA1Ufmvcf2w
Do5ZdWaguQym1BI/AmpppTfOwR3WRXGDxKHzB0hbsl7r2tZIjaYuLNsmkIGyg6PevqebuQIBqHvV
4VfTTh5Ro8Lo+HeoflC2G5ADp8VIEERmo45Qmp11svTlIpP8YIs5LWFxspamR/Lq+QRfRxd0NZaz
2AOoY1lI29jdn1vmckOJevQZkNI7T5TLNc1seMGxenWX7OefNOM20hQa1MVBl9BG0IrV9w99QiRI
Zt4mSNL0/vwoQC+/u0aKRzbHhs19/L4AXlVl9WPiBozNZEstd/h9YIJmuyj3Li7juayQZoVE/gf6
5vE5v28DXVucEDTcjMq3PmSnDjVYtLPrDuOm7XGIVef9f+Heszk5rdtS8d9SsvNJbjrNMpG21rLe
iETSuP9/109nn0uN7LfQlhxUvquZLOG7b9hiv/TXMmJfP0dOg3nJbdYIKRms7mzGPKlko3W2cyYc
Rt9q4TbAYjcn2Ngeoqwrr2xbpLXt/F9Kg28jbMFIYqtk3NNYspAnWbK28MRh0220FBbb0K42sdx/
GsxVQ7D8DBr6Zvw7EcTaZa4T0tMBv65Wa7ciNhw1MHBw/q3z/nsem+dI0wVHSp01HyY0vaNsrwWv
ljivHO3WZpJ07Vm9hJjGOdzVJeDIxVlu8fhyYtNDr5cC+Zu7Z7benWoV+JDNQKQguyXI4tz7PGmY
OEOd2S8PELZ2BWQmfOLAWNFG1O2uO2AwXfgQuNNEkBOcsDXFugN+Ek2Mp0LWrXBpvfZg7f017lvA
SfPrpaRG4w+hhb9f/kPspITlyHbNrr3bU7fO8PZb+sGTu495t92ZltdKp3jmlhffpV5ntdojI1ZU
QusaOh5ThPoelb94pWPbgQFjYFfUpfEVKKt7LBINdUNf/5P1N8P9DT0f0RYn3DgSCJelfLZNXDbi
lMw7yduWImCHUHfwjG+tGlc3iPkNIfvNm/tXRJW5v7f16DjaAxxlDv6epT19ilO1Yo/AaTX1GcAW
MQ0Gn9AS12T3idlIQCoo87OQASSNzKViFi0inFmYcv2ovJKxctbUjpNNMJtey/4r8x5zRfZke8Ri
CxeATRWZJObKHuM6+KYQ8C1TyLqdewc0iQk3wTPhtjBJhUE5sf9ylx4+Lr8Si0Fi79ufdtiWDCwi
x4Jc1T4q1PTOLhpe6FKx8a+FVRohlBOo0/o7bXKas9bCMumgQ9SGr/LWWitS/UzawwBWTIcNDj+8
CIbZv89VWZfB1cPg9MyQQt1Kyz5l0WyHSrxWW1H7LJik5fhUS8O225czBM8gmZUuzhH0g58oKrZX
4d1ZowMYbAKbURxPYB2IWZ0Pd4K05syMjL8200zlDbdA14jLoLuFCga5XXBzB88Wa/ZeoS1IJxME
vpwFKrzyJ3vHw52MLxms8/KAff65PUmozmNL9V3SgM7CYwA25ZzBd3Akx4jolg2qLypkbFlPX0TX
qd/kj1w32SFWbiEdyrO3OjCsm7LlBn9ASSpbphayw8E5SGyokt0yr3XysuMfYLaoDmpd3e5q9wEV
X0a4q56tvCi/n0k5SJxh4c1LcOtYm50XsUvMDmGtGemtxLXGZm5iuCjsput3Y5wrYpxDv2sjvDWy
uceOssUtX0wPdgHXoEknUnvkJEjISGSBafG5wZbRJVCHowr4Qtr65nYqJx9dkW5v9QoOFFqyV/hG
CJb30E886HWvo/9AwIKx/E50RKR9jB5INFnF9oyKT6q7hHBuhvnlbLV+a/GBeBFfNvA+3PR+vjR9
YDEpi+R90RzXpQ+00CW9QlWSXfkhJipr2OeaDowGK2U1GA7oVBi8AVycQ4GpFfhzJjCjKLYD9W7Z
rULlzhM3a/7dZv/+Vu+dh143SDu8NPFdlm4L+GCT19udW1TKgkdX9En2yaXVILPbSbczfw2mHoF3
/YVs2vl3X1nUwlTtoiCpqwKw60i1Gs8TbONVFTZN6hhYVDnUNw6F41+0SRqqy8OUBTWVRc/HbGIT
SgeZbpVAc5JwGVjQqRM3mP+8QpG9Ffn09gYwZD3Htr5XXxrfRP3nXsSPKSMuMTgXXoMTlJtVgwIh
PDozGGJREbANhbYg5kmnVi+/LMfzyO7hOwaJWdj8UDfjBxj3zD1okvHfVwvpu2FbISYYnHqRXiun
+6gxTae48gK9yBK2NdVB6z1e5HgcX8Pz7qIzmJLT9CyKqqPUjZMSiNY7MaxdYGrb6GU/g5gOLWm8
95ZAiKMYF6i5X+En2XDU7onZt0iqOQtQBYM9uLXgawOq5FVOxG/eG3S6YJYDk5P5o+PD9qfV7Ela
aKhnlsUY/vWjXpUhB5/jS9PWSUVSN+7vrNXTR5j+9vC3srL81fPqXReb9Q+CGSHKe6vfEf/U0wJG
44eQTcgdPuvykrjL5DmQM1TWaucTeH91qWIuTRpxYzGYanSmw9wQ3I7gAdmLDCRnHW23eC5zQUOt
Z4GqMtDTSZHP64CArp6fHxA52HjzaRun+q721WDUr2evvT5MedvRiWgo4Yh21NWc7rUAwKFZtEb5
FxMXbWSDG27EFxZ7ZAXV1VVevaAOFMVQoPdq8WjHFj6XGaHI2oJUbTBxknqqHOlr4RqP+aLLi34b
SvbjvZ7/9pFYc6bZ7oXsTBFm6qS2onu4Zp4LiLYNkrsRiZlMIfSMR4eGg597rp1bRzr0W/Tl3Lnm
IAqU5DafLBzgUKC2weaqjOXN5FMdsMKhyH2GfcB45wCuK0cn/qMvT1B96tuUuJkU7DIQBUG5LnLk
cUalWMKTsJasNjGjaeXIb4yishP35Xq8iloS1WfAzw8Pr/YVareijBXn5DL0s3h8sk18oQmQ4L3Z
FGWaI4hADEjVwSxstTH2HYa7Ni7TKvjtHxFdmA3yb1TnkSaNXroP13SewrcsZia11IxI7z4PqG7P
hg7btqX+/zgg2/F24NNmaBc/97O0xvBFg33xxve76cgQ5qf8jpufZwAy5xdH9TylD/z/XZ2pIsm6
Bm0JircfxrNMMC8/uNR2OpxoLaLR6uDEBAGDfKoJDLorwBbgH3zhP1rwy+lr6yN46Lx0a1loKmVa
MrbeZ1cS+RrLKnXQyC1kHM/0j5ndi/hih3eXgMNTlxQCZx/voVXe60+u8Ynr7Y3irX8mN2ngjAcS
Rd1mteWpvAVRRX7D0QR3FBbKrEs7cMQoSjmn8ZIl1f+QbGm3kiBCV0eOzdh/QxSAeq0coBV3dQkd
pLMg5RuoFgAFrB0ljvif0sC1hSBuwTHuRE8Ov9eiOSc9TrzmDsZJ4KXdevvoRGe+wie6us5NKSEQ
TWzqPfnsZ+eQ5EUFqmbZerH8HttpegsERMom86h8YpG00XQS0VYzMQulUzW463ey4ZhookAczLaO
45sIDvSPkduQS2i8Fus3Lkh7W36XyNM8MIHm9eZXPs8GLpnVt0a6Jk6H5qOysEQ9jn1gWDkEps22
NiWNAFODWu8qE0kf8G+fEYjq1xQCRh8WssxlkIyiQyr1YgSa/oUi5Ed3ZRXzet20CycFqDbsrbbV
uMTXOQ4Q+4AW4zqM/IrKXid8WRv5+TjFIglKLnyQI/f9qMug1P7nZuJm0LsOLwMd8DCEa9jmLwdy
vYaes6SjE34PQJgvnC9m7Aubr+IgkeKf0oZGafJXSUF6kgk0jEmshaC3yn6VgwRMD9Mj2Re5pDId
BGjrcD1Qn0ik9WFv6874g5Ody6FsDA6Ppkno5Ku2v9/WOdSQ+LNwKFhkPxctt85xnO1xeGAbNK8J
unkkzSu97OX9Tu63pIw3GDd+RM80Ym4C5Ml6T9RiR1kzpXfkHYuWEN5NV30L4eQFTZFU+1bvyO+N
VAUoRMoQp4o5ZlQSOZkjV/Bgvk4Z8AHn98BPiSSBLmaemotJcglWM9CaHAj+cEB0vDTHhIZ1B6jm
Ib7ExjLoC9I8tQimKRad6rJGzgzz1YAtFwajqPg25vTO7KyyeJPLp9pOLCcIzGozonhJoKQ13F+p
3QxWbfPeVWnjFe8ggpg5H7V+WKaA7Jmc7WBsr2YYrOFhl89ROxPhoFrd+GZh+6VYO88RwTlROpAh
wBERSnLm62r4+zPkqjwDnW3b19ut8cPLkKNNj1JEsu397KGEb+OvLqQSI7BpmBr8CNpXehPgpSx5
7Vuq5JdUG7FGyzesrwNHsxuOFLPpy4yhkjXm9EsPIlx/h5qRoq4v3cYEbFuKLhFagjwKs1IsxuXX
KcAPuQiuVcptZVMsvkkb0IitqTXdPrnGeOxUv7iRhSlja3XZNhHonice30q5HW+3u5+mou3cXf5O
S2+4XADS7eaFkqtrWJLu/gRQGMrQaKPVdO3hv1GoCUXY7/DTaSbzvL+l7bFk4DbyIbWk4Oez3oci
8sNY80iflqP9mXmpUPi/ezYY+RPHbhzdAZ7osc1jfv1EjIiyuTC3dBi7fwuDWHtnqra56drPog1+
hFei6nEMBwVOqzCgN34l2OoeBfmxQUIDrzWjIkb2wpJHG9QWwmgiyrHIVRko/ZVXp5SpuKlL6YyJ
H/Vce/tN6dxuSBlffM1FWso5wKBfyybcagzvDbvfKpfjldYnX7VAQCbKhBsBfeyGn+mpIO/maIFe
5aYBdpEmsIJfi+R1e1KJ9nAVlfORZhuysFoa/VJOC2TWlp6Ize0YRz2wQ9PZjoubNMF3PFoxjxkO
62J13WvOsSRh32Wm++FGETZPs+k37Yl1oxCyXA4QnWXZD+E8/K0W+mZdJcRuj2lhi928ovRVZIdg
UwcEY8W5e52oSwYUN0Qnsxq4x2N+SAusjKlVVclTVye8th7n5ncHG4zJ3McmP+Au1j/Tp2IxiuqE
EwqXOZPOTLd3tAZyCW63zKltD8m0oGlyDmYKgUQFKYCCYLASOQgZWkV3joXZuW9VtyZ9RFE2Rt2s
HVPBhh7Lk0iB54My73mwwSg9UWd4yE+b+on5Jmr9lDlQWKS3kjsYSFocuixLFA+N5LDeT6YT8d4a
nvhxdxrWe7fegUh6jIg+0vINu/IbF24pFcw/Y5IIt9BOXUYw8qKvinXfi24jXratysWNggFZdozi
deH2j72yS0Tj+ZZTAKRQBHRdWliVCMNpQKQJjgXQsz0PWlKm0RVzVxMOsQ+uoUySaDMMBY5WmTYp
+zQ+qE7Mku+1fNcrRgF0y1eupKhr03kROVWuOV5mNYwvbVhXK//yZL9e9owhlQX1H+uMOpuLf8UE
zphgh3NWQwoRsTKR4+pCH90I9cd4IOFwUBLLiNqgXVKlqN/hYq1Sdz6p/UM+O9Pfm7tgYg80k7I+
JNbqoM+qHDtLIx7wdN2lPWMafjXq813RjMzTtvKrFZcCP6IJ8Uds/VdCDVlY8ngzhJHpCOgnH8am
jvEuwO/wxe5gkWxSpc4s20sJcw0yMjsDVmOwy7oz65gy8aPEFpi/GVCD9ncR3EORa1+muwfiKNCY
cYWQLSZ4QXD+vQ5ATajeuWlhZILiRghFDzbZwH4+FkPzMgTxEv3hXy19BSlQ8jBBHP9lRS2qwZJI
rcsGRbYGtQy0jRLuNNXEp6twyrfWh2hHONfGpU4OtDoqBxVARE3OoyJjIGQ4HSvVgAa3LeBEwJMq
UrllXoZwoEEU6zveWC/7LEyZceDUgXEA3ZGgXO1WHGHGRB/bzZobT73BELBw0ienKHZn6e5QvegQ
qVwqntYjMQjKakAMIsUUf/vBRqydB5KCwnBvytjYM3MzeOhLmrobfTo2lJsBg71vXQOlaBoAWQos
qG8eC0Gy8slyaIvTtkNfyJz1BIcD2ojO1PxfHl8IDdXkTacvAgswHskp8xC8BR1GpUt1CrTcHeSb
QT7rpzIzIYXy+PmUbYbEMAVhlvgFqmrvAmfYZtyxRbfb8E1625g60VBNBfQDG7SNPH0bPZ0VjPfh
hXeNIuE/oxMZGo2zA7k+h3h0bTKrjgJCdGu9vA088DKEzZbXHKwDUaJM1IMCZAIBmN0U7nu/1qp8
BR68N9dZMTPD5K+BN+iLCyK3mpaV21IeYfaKMyME9b9+6piGxr3RprbBc7URayxl4aFbZ9+xhvmW
IM9ScMbA3WRYFS1hXxhVSyCbC7vOG73e/HUUIP1/gWf/yNyvu3tmqIeDozqYJ3A5hNQslgpGst7a
yYAhDr43Q/mwdTNG6Ht6igyN0MOLF5cz0xaOEl8Bo+4/xJKJAkhpd/SkjGuenECjvl2FrEePHyjl
8Dy878FY6j7jq9iMJh+KAJfBMh9TInNbAJwutJEiv5TdItYra48FMFpNawbEqu1zwRJvc5OlSrtf
O+V3S/BlZpQaulYG/wcerKhUstSaN35sX1By097szWQjhG/km9c5HEAcnEi5tIIDk0dVvmWSrwfg
7hkfNns97L7jhXlBvWHriBclDQb+4cMfWLLUd5EZR5BDuJ+59y2THU0/dYxj/PQ05zoi1Vt9o9O3
+Q2VuwYmA7TaSt+RWg5n9ChfWV5sFFhk0q2SFxZw97h6WMVPf9PD6RpYty8/EKnymdDEtoF1s9Ow
U0psx783MEzslKo9Vsz5o5PHi8hb0yirw8WRwAYRhBcErLVbcEwURVB2UK4R5YKRANNhFeUm/2W/
TeIkm1ZWkXevMnEvFSltege7MPhKrQWxSOBCYRbJRqHUxQiX/vhsVcTdsGbBAxD68XFVMOLEJLWy
tktA0yvGB3HPndfeortkr3IsGiKLN8+9KMU44PpDiydFNtnRuX674Jq9Onh6M5Z+qreiKRzjpLBe
f2muPhS4GtnhQ0l+dBipLPeLplp04ADjV3+ZoU35c+gIXMWCwRzMrJ0pnllsFKMO4QtXspt2OV82
0bpx51uVV5Xc3NNK+Pq7t/W8jLHxYgvpY4cnwUNQEWcTI+1CuGVXUVR8od4LgUVuzwZdlI5mf6t8
ZUnlGGvVT8hyeuyzq4AC6ifKWpWM/6JAukLwLRg9kmWrX7LyS/yQJWsDHXMCLAQTCbKQte0jzJm9
ti7pSFwht15ksFhGbB2EJt7T98uc8B58PxWBcDIDiGLG7hnbm5udDaIOKr2nGi9mTHe/bbhQv7jv
nYIBF8F8C6ze8cRgDLcTdxR0JVF7CQPVMbcyok2kwJD0Xy2O6z8Msb3BrOfQaxwmMLtJ4HBtmfCg
ESlO/oMPxKNHnazaaiuvZonzgYF8PbM8+XCgFH7hYvMEisGQ0mXgJ52BFqtUPrsO/T728r9kI4cB
oRQnwZkGF+Pe4mcZlSiK5e/oUrqtFAm8cJtf0c/C1IptjMWp8VEdIoA1fER5DyAxg+XBhE60ErPc
3XqBRAaTTpCY0BI3iIxI/LfrJJxU8a8KKmsJjZbZoZyCGw+p/fsOYIp1N5D6Mrv+Ayn8X4yxxjQs
ADOoKHN10fUWS5YZ8fN03Vef8HIlipnT0eh50VILpPx5GIoqw0g+r4HZMFNDyNakLZgaOB4LJgGg
SyVT9yw9PypHkrvLOym/lNf5NBhUM7mDOW0g0eiOluK3fz2Q5XRqG25g1NBzy6Dsz5XOGQ3+i4C0
SD9UUjhPZK7aR7Zbc5QbWEcrPYJHT0NZ1C0QHwQNafcdT8C2c6sViwjk3NPPbbxrQ2JmcS9M5+w1
jqkpSwxmxmKbG2e4Ylfa86X0gkflZ5BrEzCenAd8FfWqb4pM2uw1Nm1gpdwJ2rnyuj9W58DNeFhl
JOBA0hkAFlcmm8G5TC08H3F6p/ENiSAZdWG3OmGNrYsbmPtnuY31fhbgLOBeHmDPC3B0Mg72fdw/
B1m4AN2JJrnJHXUxEWV03U6z5WcHZ9fUDi3gIunmW7XRCobW1onF4220uZ9FA1LBg+C5BDq8kPyy
Ypn3kL/TORaVaojqm+yiT/zs2GxOOn7j5tV0hZpX1tNOfXMdRMDQgzB+xHor/gl4my1vZRFmhgRR
eOBiS3cAHC3/1CdSe/dsW8uBSHNCEs+Ak1CPvL8uHvLcwo8Txl7icq4MbLeDdBtbblMc1hTaIgmu
NesXfI+6oZB+DG4tjhUmf20ANSHUNYx9OrhRH4Tj0xBZRlKnEZbT64TiGLSkOC0/ZsgoAPR6+Lfc
kWTptS2gH9TDQAkpbA1C9fLx7A7KrRf4m5LbzaXlc+01Li5+8c1Zxn1EOKMdQWBOzxJx82FnA5a/
tTeZG4A+4CmH/7FV1hSF9k91ZUex6YPSWtpHAJGiip2ReBAEFrcZKeNo0qdzzb4Pd15+dV89JLYE
LecCe5zk7lIALyenb8a0JmYT+fnQgq15o0RnzerNsxDc4VHZSVcykbUEgoXFpCWy2Vt7a3SEq+rF
qkU2RWplEZxmvMw3KLVqmg6YcaoILCLPJkjbQxvSB8F0mdteohaBfVFVAp9JFvJUweORK2aTLz1I
SxmcsJxdpkpwZvB7c3860wuRb0YOJqpbwYoUd5ryhivRm2r8XuKrUZCfWUbvmVzSxFY/xq0bIaFg
0/wYed2DiLifCfIkm2gK0r7bIcfnCQDaFOecGLBQ3wxqP1pfpymp0bL1dhA8Hu7AwIykjgCsODZM
35sTAF9hkDjWu9/7kNLdrw8OLJBjHaazzcYMAIH1RbEUHculhI6OaTgtZI4vf5OJmHYnPlYAy4wm
dlKpPl47DduQHuOXnUnr2gACNnoYLtHhnDXT/3x4iJ0VoMmpSizxb0tH1OugspV8KrneTPLCi0AK
xTV5sQZvlOsbvrvLP0mWah8V6eyU16T/xQ/k8JbTVndLFSdgf80pBmxDN7gtZr6lxfGMmkaeNzVE
4YqL6QKAv4kVh4o3Xu/fst4TBHJoDbNJ1PC0Jnuy0JeAoLWuXjfC7sjhjFVdZfUCAGTAPf7j8ui7
ZqLjx0U6/EZpqraWtK7P1XSuS0S6MA59daFMM3JMOAyFO6HMWuk4FFIyJsYoFJAVVHXT64i2gB1N
P7eGLzDd4JMo+QbyZIza7EQLeh0TUq4/mvgw99AupCs/nlcTH9E6tAoOvjtXgGsl4o8Ny8uVsPyL
RzzneaeLKJbOH3tournbv20d2cOTFQnrmszj8IO5NU+ya3eenq+sGuj4nFsffiZWXCIk360s8xkV
hsnhkZw7Qj48vWy3nZhkzKMc+yeofFQQ3LzNqHeJMP7SEG0TJ/ZVVfoKeAzO2tBIBqWxyOVLfcm0
XF6lggafB6YC87JRG0zMp/nx/2UUAGNFVJTb7bq3Aqksrb1MdgBH22PTq4wZ2g1OIiTVgZhQTDx4
n8bB7WigPWH0NkmB3VurqIcGcoi9zPovBuuByzD7MNNyromohFOFDECNwFEGdwbOE2EvykwNRzY+
eMirgbU6LeH1ySlLsxIIeP+KkL7xuJjtFRh4cNXPPlxdnD0NXlFznpT/qKGDEIpunTuXfnXdpnvw
NZE5bhB0vHrpeA6Ngn7s/iTlKJSRtY9R+2mpWvTGbP/F/ykrmvEDpZo9EprNalSXJSoDJC5NmiES
nlc3nIteK0JOwOBXtXqO2gq/6fmUNxf9hE4tMm8CpbSUbuoPGRZ57j0tgGcYwvppjx678ZwEjRJi
tx8eLGUk9bKh+9LmDQhd7NFDmgKlBIYE/MQsYvw2WnnsJz/XGzlz4qQw/tS66eSBwya+8SvZivFJ
HkOgoQWTqZjFiGqJ9IgC8s29ZLDgEf857/JUauqu+rmcuSqv43JQmfqs9hxAIH8u02NbGOGXBJLc
3/5Y9xv+2hCQIwmIHa/gQZRcBpQKRHTAIUGR5iA1NLPdrfz74x0Ga6rMLI/iNZZmKdylZEN9TAKF
PdIBjq4UkU8vryPB6dq1ImTQ36gcQqA3cafyj1PcNEjkH8GiVuLNfsC6uepw+ybfpkNE9Gr+x8cb
ikt1xTUn9jz0YbHB5+QNA64aeaYKKiKHHmgqry/pjg8gxCJgAIikDVo7a0DqfIoCvhCBI1IWiklP
DbGWuzcIPF6D4ctvvVL7pMt95D/7NuF0Ueuc/qe+0vSua9zb7kTPn+ROEDDDzbceU6C6BgrTH3CU
DaRmKzK9y8ddGQ+G17hyx39GEUWP3N0TL8sOpzpFVXgQqXb4QMmgIwT7NL8sS6egBDRBb57E8nCy
JQLSusUG0q7K92iC9CkQtI6MY5nhgsSmdRMUmvROyJImNWzTrV4nL0BI3pkx+jLGqXSUyWnU9Bl5
n6hEy9booXe7MgL6gI6S1XIQZqhVLIax7+F2Wz4zJn9VUFc6FHnxTyoJjxebdOvw92t2BYGnU4YF
yHJLLYJrgAw1uL1vYrmB516FDODisIXRGiJt/EjVlsEjkT2H+0d2c93AvTo3l9zT4yp/nqSDTJjN
o3zhXm4omIfa32SmzFVojJQ+NGqoR/QTUXQTyfdDA+dZ8tqH1pSipHuUEaAJDM7MXdgBoozUfjBU
Fne+XzR6izGfip/Psxs3t1np4OcjcF4uMTgtdKovtwYEEICZfx0I8FkvPGiMm3CMa2it/B0CkBJ8
665ktqPPe71Fsk9zf4qEkdXuJZ1NmlFD3NbVYCCEJYr5il87dutQaTOjuBlJ51jDCDH+X8EaJFqT
Pmf6mleAod2w3Ve0/axFRPyHDdhKjrDCfIt0RxKBsBVSRF+vuonNUUe1CesHNrEEtnjgu/VOIJEp
DgIzGz497Zwl3Uni62iqIPDYjKvwiDObc329m/v6HQ7zrDF7XGRSiH+m7ZpYgFevDiuU9cjkogMM
Lb4jHopUf3IypVB3cNSO3QeUCj1bGhvt1UKRi0m1Dkoo/he3IlsXVqR6hZ9Rw9hQwLCu1jtCmb2c
fhFLbrdh56a4jq/BeGBSgt1Amr5uFdjAykm2KPM+eacCKowcB8CTpKmP2s+X7FDDPga0zJVCwSYs
vB+KrQvbu3kRNhn6YAb5raP1NxNWpuQVcGmELDa+BYvRzD6ooSq6Miuf03GljaS2QNAluiyY1Lj/
bg9mwkYOmTqegDGFk2qA/ImP5MeuIKAGJM3jPsmKBnIe7bPjctXssa9TY6oVXZMqwOWcyCVTXwKL
vRIh8EKW2UnpzjwqHWi98dyYY6Z9gaG6DQewmplC7A/q2psrCs7OwgapdLBFeHXk/BJqvKUfPOGf
6fWKtwPrTMFEbYcQ3JChbaGBv2hVmJbraVrpVNFwXCaA2FZgC4WQVmUZo+MGjcgRwc6qSz8TgUEg
1DDuMwkiIXQ5QKdJhq/I9ktOyxEBoksNHaxwmIlzd2cXUuQkY6fagePtZ9IaijVf2QPP/IkH9Uei
0apYM1lmMOI+nWy26e8d5DTzNAhaMjuYe2Ao7Uja9EaisGH92xzFCy5pMD6LUuGT1vpR9+h8iOYX
1ZiMHOWzNZ+V4p10/cr614/yKfYG/Bx4mbnebBY4MfRW/pI6alsMCS9mfas07frXUmcqkj4nVJI2
wO9XNd+SeDNJ7M6ZWVuomoUM/zgw7tC/rtYXz0CE2E1vD6u5hMtBEVeauGXPo3zmvkNfyBuPvfSS
dO50msgrKWitX0t3GLRhVxmMmH7dH8cASEo7joUxgiyxVrUD7UADdoKkz7GlXwwEij0A8/69CW4g
SjGDd4n/I9zAFtWyqSiAV4myRKwGQwswi+gUQuEfirX1j7uw1tzIOpH2bElbn6A5XDXhkt3FROMV
PXRDLxS6RjCu5NOtaWN4tgaRCvCcjBFlBdYTZC0R1U4E8iOMMNZbMTx9ewBVl4zbzZu80z55JNGi
SGjQ/pW8pZ4+b/Uxh3ra1CfQTa2Phy2gqdOTWcL/9OqB8MCcyF9NmnKexabmDwL8FkkFaAnF1Op3
64CzMLpXxz+eGz0HqakKI6eFafIOQDOgbaH1L2N5soAXdQZK8BeSrW2HTmjS8q4GvVzrJIKVsLbw
wLQl+Sdm0nHlxNF/K9jAg2fWesJawQbBKONOX34TLj2HTuHzewQIBn3ph211POimaSBfcOqW9CN9
dg1Tt+oitXwe53qNw6sl1wpjjdPyprkVow01VzWX8Kt834JajwkmvoTe2TO2/4sq3IWvyUqHv+yN
eNUTY1ZS57ytJ7EBx2gdPbHdpag+LBpHJcVKzgT33M8cq/vZeoItZMEeNVWuWsh2iMKy7coESeW5
3Fm6lknxFHUqw5oQwuxa36xTLNcsffgsQSA31VL3RywyHDaafWz+JUV4wDQnHsyf9rWY00I9/X88
umTx+hiiF7n9arWbh0vTIHwPTs5afYXy8nuILVVedKPsF8wQTAu8VZWLE1fIte/wukUNiBkHO78m
rp/vmLCrOY4NwgEzYI3VI+nvPmVWfdKuhR9cjw08PVOqopwmtiBKMDsXyUix3+LPwzvBjMZoCiI4
3m2mGZPgqXqULnwl20eAEs36dhNBTJhl1dpDRrl648OyVgyOEZXj4XqKn2Q5JpA2nSiem4jEKhe7
RkaKS0QtOBr4qFKTs23jEkANZ9hyLDuB4Vtrgl2O6iECoHh8elrcLg4QVvAkz7tVRYnnChSG+ij1
TVPJsk5M9lUc6SF9tY6A2gtxXupxlLWzdzsyZ/LEHK8DuSbuOvrMSI0z4V5i2U6fcmMlcpMGPYyX
8QRVXdRnPMeVoprZWoiy3k8bV7pjF1pTCMGC/NuZ7p4OqSKipn0XCwjwiHvxscg90x/Y3fbHyJuK
MUm8kn/DeBFtT1DVzhoOhBTvUsvGrwaOSk0I4BrF00O9ujqt+1ocjjrRm757eOaeuKiVqN482z44
najFHS1Q0d8U2q0P3uZp6hmN5+XNLSI+29bhHY9vjAfBVN/6YW3aQ5NKZ2FAhOwBC4z3lYvHyC+d
b647ZMNQlIX7T9gOenmZk/Er/xBeFI6d5x9zV0SdOsfiLTvZyY58mAWtfaUY61P3DjmuKRVSiTHN
nPl4EpLdiE0nN4oJu0wg+kg/KbZVcx5khzp6plcqYCzNt4Rnkrzj39JE+8iHNJtbTHbOJuhYHmBa
XBCPeL5r/mFrpfpyrT34dxrVDa1usSZkymgNh/UEzKSgx83AfjAVdU02mZ82z7gZuQOaoHRnzggm
8thYFxOcvBo+86KHKelavreuAGDw1Ya3gJHTjRETRgnQPsfcPOC7yHY4LqAlm3GD/BhvSoWgDlYZ
uG//K9cEgTVGa4QELDRFZsbtRs2aeLm+VT8KoDagQFqQczE5ETvR6OuEhw7F6/zQxFnpRnSZYXyc
G6hYeNL9TNPV6HkIxwOIrvRQuTvxLM3lTBTTrSgGAFBViNvU0NQ8uLHT4zmLjHZJAvWLYedMi0B0
wJCUtWEfmFoeT8/gG04SWcnC1j857BSlkw3ldBaoSM5p9bh0i5+iFMnvuOwzTdbJgUWCIi1iQyr+
vnvw1v9cRIDW3IY2hoMzvRifgI273nWsY4oFfvw3Cqa/AxKbQfmMOuweworsCxUu0fFwon8NKS4v
kzTTfosXBzRQIFu1OpJlJGjcgtelTNJEjmt2R1c/YAwJX9cQ3wWAbnALLGEfvI9yPvGbKfmHXn1U
g4FYxb7MwBte/LPJY7Zlge6k5suxY4+mddtRwPNMItKRydaiixhO3lnHBnZP9nLlvZmTGwO1D+55
fRDQ/Nl8oVF04/Vo2CCD1jDIUQGNSnCIYHrGjTrT6MmXkXeF40nV08tFquoK1YVk5KNne8ba9ZWc
lhwTBkJvO+DnZIhylC72I5HgurGaczEZOQI5ExBlqg+Wdo+GMDJeJTBbSg0V5pQG18hgXejLfycO
YPd07DZ7axohijM3wUZd9WMGQWL2ldA0XN/Yj/nexY7G4YKYs1x40hY572ncuN73dvvVZboThZWG
h3L7TddieAV2TKm2cQQA8UuihwSCWwujBVqAMCBP4wFI/ojMnmntuaR6WdqRSb0fvmwoAa3cPt++
/mA+mbp+mWB6bmKYK0zuXjGRV5HlX+FXEyxZJMZK2FA70N64EeY746dqDGbtHDdro21cyh851u70
YwCXy4U9ojUAH/v73vwYG8AXOVRyAcPdUqQb+KXE0PIVqiBGpw48I+y+vYEp4BtX7jdF9tdyArJD
tBo0w7j452q140lyICUdXIqYAD3HqFJIsSvAT1OiyN5/XBVeT+WSmN5tXEwvf/FyifL2N2XPen6u
uFCADtfxkdzIx0TseRD25aAEHAQ4Sls2aOXATWLLvkTIerM2jLwFjKY+u8unc4pwPCKyNbca6SRY
h/PH6NYKlhxfvisksjtjsXhdkB3t/oiQ9dSo5JcXb5uiWQkr3GRUUdbKL7bu7K2uGbzuj5J/2cRb
0dfn2AaT5x/nRRIAUUdJrY3GyC6PmGU+W0dCH4VnBKKIj5Y1YrPbxGvIgOyS34Rmy4T0u8mxVM25
dPj/xdzCB85F0Dm/ZANvs7+GLrM2WzO8Q9cnxrpuQ9tNbh6HO1okXvVNETOaAeGKE4fiMRck0uix
xbUqaJx9kR6xSeCS8lISJvQtkTAlmiUE7XpiAlTfqrMjHu48IWqGzBcvMAMXHf8BKBJ2Hl8FdPTJ
a4YddZmzri7E41lh3NaI5WtbQDZW+H3pvmAaaiLMIzY38Gv044AKZYxk34KHP2vfuJTfacOVtCff
7I9p1ocndU889nCx5OJwejcKE9FA7829vpfv4o3opLyFgirYdcbC3VmSO67TGrn06VmfUvQ6Iv5c
G2ajVTS1boG9871lQz60T8WkBOJX3UphQv8yU8UMD0mvLNvMXY49IwbcJnVtwppzlj97XLkoOrPP
HEZ5/5XwhWSFkEuaHTNiKF3WNoAbVbamK4EIjwK7avMvAO9Y9IFBvSKjEWk0+8PwPC5AP3wzOpuR
E7TBLJhDUHyylJuLLTY0aIZs/8/0fObsS4At7gGqR5NDz35u6D/VWInB+Cp6wI9aDFhm7bw9CTfw
DX85J7pGabh04Y5IKRiMUprwlPJQDvOhd1MR5sReCT3TR9Z6N/gSUFKMykU/M0SpQBSABQz6gQLr
Fis2MdZ9OAvxDYDt4zgBhZ56/j2bGAwnFXBNygujUhK13nMssdDbIrTW1qkMFy1BgaEvo5Qvr4GN
h2l7b2tA6KN4O1/B61PzEu//3avvJiYbTM4VlOpFmjG+3PTY5J/k/Fs+IvCq1xjS8CvNIaRIPi0z
DT7B7Tkbfl6DG+NDQxA1bNQDQcTaPjPRgCcM65EUPCj47wm4HiWC4jwKLwfg8YIRloNqMlGTw/e5
iKoHxx4bM3TgnARUPipMxoSjlvZp8W/mUr5wTlgzuzOyhcxVBHopBX6uapwREQOo0lmWN3EZZYhl
P036zkP4OLeubXWS9QTmpYvq93C5KJ/IV210t8Pv7nRvTuTMSSoYThJ97roDCABfha4nCm1R8Woq
QtmyPhM6AWVjZBsX2hkHyjHugZ//flbM99DU7eRBcYnHr6+j7nUT7eYsAl5e5enOVV4n1yT5VOJr
wC67hQGVsto/XPhBra6CAR1FM+d+gfLprC59AfcvcokA4Y0qDCWrFFg/36pU17guVnxgGD3ROnxe
EGlr/YsRJAt7XSYM8nq9x6MtqFhkhbFi1+xqDr7b882uZpq4ME3yVaSVC0iGrgPrBxVhf5HTdzVw
UluIg1fk4fvhmKOhrBXbEMGiKipuxGu/4cc2W4BJFcFNG4iGehYi08Mnf6oTJmvevtCOGvfngJr5
HtyQAJ/P1aV5fIWvj9WnKGWT3OUiDQxJ9AjM4pUXRlpKjjV/8QO+4skRwpy7j0MHAbP5E4QO4Onu
scyME4i06XFsufu6rRQIP7Rmt1hLDtpdsd33Vq/rzUrvWBli/KlOe44i5YzcJ9+bKP1GTVc5+CGr
p2gqdSd5J5Tfr5FJ0fP2ZpmrxYm8lIZu+z6X4/mr48uhR/6KKw8xwX1P5FfdOcIdPRFBMuNlofd4
Q3pzYQ6TaJzfRAZRjpV6tG6PmYUVLYdmIUJOBC3pZCmsrOt7ehd5kCjghM5tFiSOImQZ6qV6nUYU
+iDt7tif04FBNodzBt/v0Nq62dlwCXbFXOgqQwCRj/wbEbWiF6U6sk3jeu83OtVebsdw1dofwExI
T4Hdjin/HGj6NICyeyUZqdSt+WQkN0xfcWQcr+Vqx+zzIsPvXVjhA43ctned5oLRf83vr6hc05H0
OGD6IZyjLN4sD22u60eyJj3qrmn15/imGGplSSp4lvSkHdBrURvRZXvvhmgiNGdXCtrWEYZD9UI1
qXHsopARkhPLZ47TiwSS4X2ENuytROKlu5RmY1fwT7sHFdl1hlKCG3o8XseyNgqNVwt2aCmdirRT
bg+KWd5YE2F+RXxzuvPgO+A8neuQvGYUXtw+raUKn5lbAhk/Bk+F/pkWmLa4Fv/VtR/c9MbV2kvI
FtnFafw7osmGTMvN8a9zV8S7v3Dbv5T3tv4rFdgqLNTj1dvCtneCxKLjVWJmOZSmP6DfTeycvI1m
LnVG0Rgqe0cIm/DLmKad3XcHZPJOxkuxhxkXtcGBjLMFTnnrexBDR5cxWkC+9hiHvBqTkgJ88+X6
8M3rgilmG/cSfAl5eKfTOCoqEWJfzQ0EhlTgcvI66FAJJeeTHsSWXT+u81NDRJu/VXGEFTJInHIl
gIXVCxSr+2o20ofe9i4xqo5dBTp5py+ODUJhVgupB7tVfEWHhf8BFWGvFt+eY7qschGBTfy1iyEm
F5+ljxQs8NbmkDo1jEy/NkRTK6STI6KKhNrTvhWAvNRN84jtjCemGa51WbEr4PxsZTsYg3kuzfXk
mMe7R5KA7aZf0HLD4RC3vn2zGdd9w3m/H1dea7p/kpD5mbMp9MrFcmD7zyDsPNB9hH28yAs1Lj5e
sLkVp2pmONbVOLOq3tYeKnJBcehWe+WumkH24frWGCXC+00KJhL/g07ijKW39v+ZQbsjWihuRP62
8NqVWITwMWi7ZEuEStY6trdZ7edR3kGAiD/kvw7eu4sBg990LkNusmoS/lUk9TV5MT52FNjTnhjT
ei/zpF/ZW/Hl8kJRTiisWL8WWxFRUUJERAMcWEHRFomxyvIEiSe+xasxNCT/DVMVCuMhQ190U/MX
mlLiZHNFYWxhq+/6xqmVEnl60LNSoTkhgVvZcwCvpA6cxGwMiJyYCJnlMW7WTwRH9W0CZWH4448Y
BlQeoPeJ8WUZn98oq1X6KfiJrImG5JfMkA84as+rqceqa/61PibimspRw1i92/HSrKonuYhynZK0
dfZpLQwzQmxBy8Gwiy5v4BN7yr56IU08sYrTI9Mb+vph4DiPbIT8z16tl/vMmD6+I5KiLAboaFeJ
mONiwOPbkM7OzFXWqyNq/cPTulF0hh0erwmWhPs2qwrqsU5RdGp4sEfwpEAT0AriYEh2Yc04lcVS
m85hB3zKHnjTRhmI01F1BJfm/QHfTqgd5hfbVZQgJEyfcTAQ4F9bPgkyDWfRuFnWB2pgKeoDSzv9
Dqin+mqPO0IsWj/BFEaEavo1wuzTI3h6HEV+/1GksrUBHuBO3M+qIvO5OvIqHjQ4Hv44a5yIVx/a
rslEpR8eUIZea0yWrgPnm34GxqrEpYwyuIHNLMQiQrLjrgZEuXM1LSpPQJpAbCn/f9N1Jxj4ufa6
BtFhzKLW+LHAEF0WGOfVrHwUA72xYiRGHgM/Zr5GGfle89CSQAF3IeIcnHvlwSbZGF4DtQ/pJ6oS
YnI2H+pd4ku3rDzAABws0PFeST1FGxrhjgrILFxITU1mX2P6TusK+bQ++DZ9b1+3ClLx3ROJD8Ne
r6WoCjA6gu1+U7Ija86Orh+ozc5wKSIdWDRS/hXZgmqr7QCff9NvAzQ1Cm5rykcKuS7nR0lIm4ZJ
gwlxFd1meLyzO/mNq9juf0zNtQdBZJ1NeQZIDqiVgEuKJUGGs38/SjTqd/5RMJ4nCIwzwRmjkk4T
FiScsgOCnxdIk7Mz5cEPKLAAGgwjWfx8QHQ/89Bqf3itMY5HJhYs56MV5MLzOdDMcmgPM8Zh2HFV
B4m6U0QrTyb2iMSODx7xMuiGTsjDbypotheug6kREcksG3rdtcXFowL6hokNvQBrqYw01VZnoT5Y
QhdAyrwa4IMh6brM4GBFE1Kx+kXqZs7cUenXMSLsz3G7ZQCf2IJVx6nkja8KYl5w5jGMSF8KlsuB
hBafHEcFKIPEPQssRL7G6GEV/QKYO9Yr6njKoep7GEAJRy8NgNDPBqG5c834XjNCgadf8DmnCZ/J
86VayhkmJzooyNNYHKwaCIgEpn1GLmkuRUtsrJ/zsRgCDhQZCwVqT3W6V9jn7gubm5Q0E1GgMsai
FyYAPpekfrCYmG05u3wrbzyG4qa6lBME21tJA3vwXejSGAsHyCcdoRsc8NuyH1GqbHEW9hS3MFOS
3s5XvRNra//Gke5vnZQOoWJWChbtJlTHU83qDgyToOmsfpaGY1khiMQ1gjbQ3tN5ER4SWkXBQfxQ
tmil5U45MIKtQtSOBK0xsmfwvDuzopL7x0deEm0Q1wyTFCijc3zVq+P/9tJlfgOM6QM55TycguF7
iFqW7k6M63fAnOuvgC8AEt0JgI1qA4AmS0HVvQ8McLM+9s3BxGr4yrqnS47zcxD96aW862mztgv1
sF6ZjsX0nSl1BK1dohdZYW4wttnzVibrdR8nMaMiLt0yBe9XXLGj8S++ujJNq2geiXWvuVetP9u4
rVAYrX/wF5nx+h+3q9PiNEIvtA4y5IhkSt8vq4rYbFUah6pmyy9wwHGFEwpqXb56Cr/7bpxXiHK3
TPE9LqSwYRVKTnb9RTQmvsAa0fnSKG6yJr7o4wAdLBalMJ1VsC0ZeI10nkJp4d1NA13fsB3UzxPf
i5wR8L81N0v5zGhCWlQ1hE7a9RFq5WCYbonn0pT1tRhkkc+B6yFy9LxT8HdNC+NWD2LrjUDc9bha
WOvKHdQzOSnBPHRkswL1KuclxcVq/PKGvwSQN/pEZoJGY2vZiX4Nt6SPuXRyiYsPYTaL4BTLfomK
eEscT/h6KsEusyu9O++p1YIiqZaIdGJYo9UGxG5eMNAWOHbrN3jedevgqsQO9e3fP2KTInEXRTZ/
qrn2onluYw1UjBWZwZzWmyUISi67JvvMeyskX15g+9bNqtvjx6MW6mVw6lY2USd91Eu2nOAXm2rA
4b/hIyTSuUrwdsWsWGMJNAZ11+aoOJ5YjbTcbvObIM2M0INKeKrxT23z9pDgt5QNEr7vvsrCAfKy
zPfTWRzJR59Aij9DyXrrio50p1N3FXZKBF4OG9k0gl9r9COxqv2+dAxKOcp8fL/EWGssGm0SQXpP
eT33ZIejw4yRYqr6Fvud4vJQ+kBx+kU+/OTOHw7Dlq/sdx76Pc8xaA2jbx2QqKSwDvObPB9TmrM6
jG1ttN46HdAeubO9W2/SOlamXKIEN9miDDfFtcZrKy1z6ZUB/ZpQzryg0/FXb4lbPydmYyKhF5mQ
JP1pD39vV7aK+JhcKKYigEPawzBEwHVp5oCUyQD4UpREfMw4Zz91xUDaTO9FCS3/bcVqv+YNbujH
OJpKz71K+zWHYtbFxZI9LPuf5TGkcmwipVUZ0mgSsWQ9sIVTXEXHF/KtLNM8VzUotS0C64ON9hEO
39Rx1dYvLaHsCbCYD3VMm7GUNwMcveoiSl726YgsDP5A1C1SpKf21n2HGqWBP6epyND31PtpAFmC
Aab5fLFelaTgSFb0c7KzVwcrCTMiDfbtpkVn5ksbBYRbn6A8FyGG6uRL31pE4XPB09B9/Z/32RCm
rRaP2DRaHcxKfn/gRX90yjC8QgIpzerx4XF7PQjbXXtSElqitxjOPMgHbWFOnrrJbjOkBk8SZkqu
sGg1NOrg8+cFcVDjafS6xfvGwy1KAwafvAiDzuI+oHS0hqDqCjbVNsbU063xjevRJhI+T1ILX/a4
veRSewwrQHkkydAXQI3PXl2LulWB/iir9vL8ihRSDE4xL6SXjdXKoKR/+6MwCu/XBjmD8Mwnt663
v0oV5AuaN2u8p5kMrT9ftXp2H8s6fGJF1VK2Wg8VZeSMp3Towk7hk6KexvBKCtUiRmc+gxTOmZUG
ENqEMqqmYnRLWeqUdRnH7wlHSJ1JcK5hOT3YUhP5S8IK051mA1xRUONkaOWK3S3yFGmYjNQ3dRQe
r7Gsp2YLYt7Wv+eYjDDQVkV6wkTbnUhEI0Q0kIY30e+3A6R6kG6r5mM8+H3VVILahhzcbs19Fb7c
19wjtz6RRmrPoJ80giXfG2QMdTflu3/GXiOE4bipHxmMAPzQYMThSfOSCvabc/O+K/7o9P3N8emj
IHK5EtluleWzE89l6K8w/JdCWtx0E5ABZ5yiHzIhDAeLFvDZ3MGg0PBUluD9hraOxPRUOGlVQVh4
tp/ghTyti9EiJj/TMgIEz0/uVsjY+vj0/X/nfWstx3WgZeSs29enaB79n9Ffp44ljjtcJLBRh9yn
jiMHVOv95ky+ElOHjCu/+bLXySZbh6553EV68QPnuJ3ooFY1euWxI1BxBumi4CPA81d8rnX6vZ/p
ZzsBhxLuvWdKCo8o7lGILI3AcWLbtMhksmwTJ+i75HMdyo/oTS/HnoldPCqIdvWHFxGmyYzHsZ9v
FlLHsyNkX/GEa7NpoouONpgoDZLH6mfyMs5z0yVHxYDaZFE3LP+LBNo0YUNoH6GRxmHmDDquecbH
z9mkO73zUONicfKlOatBDE+16abvkkFpG6G8Fqt0e2HjnLrmEUwVwB1tsTsAXJnNpeNgHp9UFQ1V
ZOWuNI+n9H45+Q2x6xA/0vk6KV5r9CRmR1Ri9ZgI88ruZmrVf0l0Vp6dgX9H1yJSJHTiqYA5l3Mz
Z6Pmi04OYZMm/F7it3TzvHmPYOGGd9pqUg9/JDm8kbMtyvL9h3IGDEe4JKPhJxpUHfhTynSEIq5b
9P95XNwoV7e2inl9AyA2SNSgRKUolYKZE5b7G2fRV4P/QWf57pWnnfhVhpbUhwXz+H1hmJMnxsza
GCGQCe8/KU1uljI6biijQ0SjuaBv3y+uy6+xfBh3VXA5iLq+2CLXrWbNYN5pv/K0L87PIUt78AFD
9oGBIuGmvnXNvsBGdwfsIBbeBUkECdYHMUNDbneSHJFJoYhgZ19HrCYW/rb6VnxSBiBL4LFa/LTq
Q6HeLseJIu3nsT6HqwVcu7mdU6oIyZ5pRdApd1Cn9kZTr/gZYP+h4tfZ82mGR3lH2EWMEGLPsGZi
H3czQVNLtxbTsCcWKd9twLJfLoPiOfQZFhoEcZR1p+3rn7nE380HlxyeVQ9pjM2jpvbJw4+RivqH
OpaIvy8w+5KaUdn+1ZzJp3YHlIADZyjlEn/Njhffle7EtXVbDD1Co83fxcJipD4yM5tcvZ5dNXkF
fVsHT340sEDReHN/cs1rSiuiX6Qm0L5mODP1rtZ+/xDgryUtPLJbVNeAbZkjwNI8ScuHYPVFECXl
B0pTsuhi9Gj+e1JcO++0fWNCGYwPsHRVXGZ356Bje4mieFXAm1XiacH1skZHh6GWZtpY2OLRJvqz
7BSYomD0HytctYUE18HxSu8Xx5EXZC7zmyOWXOzf2nB7lByC6HkBlIEb/x+JqSe/Vqyr6EeWuh75
Q59znykPn5zlJ/LtsiksftQ1S5I3IHSvn6y40kIaAOjwpGkrAO8E8dkbPMMTZHc8Z8Vt41vy2HLd
P+f5ueVlZHltBi4pzH18oBGqgncYQSWA/tjIyrplRDUDoa/EoWQCPDw23iHczx04GOkOue+gEHpS
0UQap/B0X7yOulfnoGAcUZ3jC2yrkJXKFgPrXQR3CewtCnGeyO5zXYUOFYgQ7LWEbYvMf5lW8AQc
82e316tf6ElR1h2+RV155nuPVWs3qhQrfY6VmzUhRPzxXdkpdkrxLW76roafT0QVlxxe6ekgmwKb
+FfglF8KypBjynzXX9OkF/mtbh3O5qECt+Wz/sFheQY0B7njRo714WAuK18VV12StshJJjJHpGQa
vXyWq5VFyE1gC5OTkYwFOOfMqe7QwO4i+/jUUTb1u2Te+ticy3y9VEbX5hf4UoCm/qu+qOtsASFi
blSDzafcYj6r790mo2+daOhFkAiNsfeeoRehjP7ICjGRrdpZbsyHhbTLds9JC+W55cpcegPX09Rj
eML8hXlGE/t3XSiWX6/V18bHqauR0jPWEyyEYgcSZY4ZoyIkvQzM9D4mTV2co+bI/J7qXaMv+X6Z
GItAcDvM5YtbOfYLXfZ5z7v4pfS1OnXh9o3CuCP/hgIuqvwWN22n6mbxMhU8Re5zfkV06B/d7rZD
4xhG0iuaxlP4/HQitkQCaUmnlVjcdaTYN7RExr6jyBDyrFU4zgF+1CqXLg2EEhlELOPzy9KDw3lr
VVoIAKT4fI6zatxXyPYHPo+AfoP/fNjQ65Al5qQV8Pv9TmZYmVRvNZs9jk2Fann6whcGLweh9FgO
rIDvzZd9rInsx8dEWX90iYJDxVQbGR7ojUt9X0O7DVAQNUFA40iulTexdEi9yw5wianDD+CHgdJL
LZf/OKDFk9+ujIqkxuEEo4knTssj7dWLjfxnVqeEbP/l5+fTAKcM0ZA7CF8TNy1rV71f+KoC0mIC
XH3FcRTctw5p1vHXAgqKBlF32mazq/0RT/tM80FI0cFL0XLFvz3zL12+MBZHBHWFZ3qXzNjs8CRR
zlGGNe/Uz2yXJC7LWWauY9RVT/7O7jSsywD80e/1oBfr6F/MiH/ngQTva2FDI968584F8r60AUu0
1MK7iayiyQTGYtZu8klGSiM5v8Kb/xH5sWCvih+k5CJWLWz4p5czrb6uRbXyNnZhWlcEzL55619L
zT33LH5JJ6nXwxv1nXYEnYP1icrmPMnYp+bjd5KQ8g+Sxj49CmUvxWQsAn1CJpxYRmsBk4LhMj2K
Tj+/8I4C95Z99SopCqadrgpIIhKHZikf0Sp2eY7WtVCmYoJFycRS+HgllThx1fdZp10UnQx2e5V9
ZUtKcmXMSQzCjPHgnNeiwufGkTWu3fAmCq2N85Ut7Kc3kChG22uHv5+nKeUBRjbA9uK/DZuHwk8g
HlfhflMxW+FGRf0P6Uml3JvAg0vnekGN1tPxWFLcvHY94HT8RymO9GmRJ2dgreYXhY33Ty1AtmlQ
4PZT+6jK4bFgJNXPkhFzLer/wufQyAA5qJT8cvOcHTqrYnxG6jJL2Ep1/IGUZipfgePYTw9hwn/H
5Nfg4LGVilBBdQlcb6VQQAI1NMe2CaykBGKaEmTj+57q2cNE2a/qcPl0fnMXjTetnyU1S+q4sOfb
B6hNm0f2gKgj5tLk2S3l8xWxUhWLBDRy4m/OvJA/0r8jSjYKXawy/2JOlB1NEqDSZg9FT19QVDUu
oCbLr6X8N2qP77NqIdU1auBBjKI1zZQ4l4auTdqa4lPNpYhpe1hw2lxtOEzVq4Qryk4wuwulFaK2
pfeNYRbbIzfgFheiwCz6XWbE4pGS1v6q0MjScrpg/8Gc75ugmqgRQlffq1TxCw8bGlClhFHGy9pc
SWFDES6wylVDMt2u1LMStfDlWnBsRG7Abu1PSH9FXzpFfA6cbWFDAKwgHFCiFgyfWrz7T2iwKD9c
AJfNIT1WCAsOkSWSaVcQn5Maboa4jtNGVG4bfnIX2VxIlr8ha1mQx2m/auo9j8+QSXZf1lHW/l0I
HMZPYver3T6qy1NrwPzFyBqQ0qWH+HMkaKBNu/qYzJsPdOT8XNd6ykPfOwCKBltPLmzaS4nzlj15
g/bGAYOrVQT5BT7ya7SOYl+eEophKIETico0n4P6QX4aGqN/9CHB27goSCIpDpyxDY9s1FG955T8
irf/O8ofeZqL3eV2GxcX9erBP2m1/qRbz/9bXu3Qoq5tPU30NTAG+219/Qly4i85uKPPWVLVh7Wj
O/MHZq1Xc0OP2JqdMVQv6TTkSM06wHKyL2CXwkbNBUDAayzGUXKf4LwrVFlywpCrkR/zIcXaLccF
GB+nHXK67TJVFDIaKBFWXUChagOS3F9rm2a6JtjZAvylPhoMVkrVqbodk1liie29aBPvSmcNeuyd
ntNjda6E2VD/6Mp0pJksQKVWxm6H3z4vL7X1NEm6/WKsRXSRgtowJoG+i/2euYfbc64awmA+XsEm
Grzy3mvnwYm945cEs/pQwPrSKnpwMoipeejSzlRS0ZzaXNGerMC4piNUYqHJaslaHE1HKFC2HSoU
Ht4nUJBszUmgfY3SnhiwFWtAULRTD5F5NckSxMA0iKjcJpT7eXlPfXN8Sk4/0FI4i09adRFsxw88
vGs1lXR1jdIgyUNZIqWo5CCLM7ZLEKfLIkcXlrQZNj24Fg8Db3I9nN0bBaLUvWYwtKM6kHtsPGDc
kE20dUtZ63QRvUGaIHPP5u+oy9TqpF/61ZbmEVza0hCLa07sIdwXMoE0dIYLXm4oGZgnITJiHs/u
ZNldup8MK57y7tnDYayjpf/xQF0kmYUmPxW4e2grCElrYkStbHWrsuuuFf8GNew2LvlpvMfj163C
2B/0UhMKOsAQOKvEPR2LthPt9xfPkyXa++rqYW+Cy7z5MSpNP4b2aavB3AFOXESwGWWp1ku9Y0qw
kLi+MvtWDIKO1n4966LmvHHGxyUje0A8kK54VJnuqO+/Po6ioK6kd/IJ6f4lqzA2xI4P2iZk7TyG
UA8tT+J46DW8pDtbfabNH/PX9YaY19rGINuW8rpcrkBNLEGQp3DkI3lx+cNuy5rorVJWjibOi+/B
31Egox3RudmkeVftcFX3MeU0xaA4wlOeXxx7X0dJbOsLMD2VAfLQcnpu3vFF1FLEbs8OjuRWz2jk
z+CVHTC+3AHiEmLnMIrS2MaYvcLjSQQ0YuDRywUI2BGAVx1M95jyBWHLp8LWdNbH38B5vnnekR5T
gd97Cdfnaj9UjRgL8a9URv1JMcLBBQd9qD6LWWKsdzAAzI6kT1XTRqGeaxP3gHIN0tR+9bRuXpn9
MnqTTi/9IzEPVSIZFh/55n+lYMSRFrRabMXZYD1fdy3/8fDB5yuOoLMepzBllUwqdbrkdGyP1UM0
7vE6qxYuLKn7NHRRz6n4Mn0s52F9tNWTnUjS7iIQbj3Jcy54sr6MLRpjtEOSkqOoSeC9+BMUsW8p
CDzpKviVDYehSD27UXOMOY1WjsqPC4d+s14fInF6WcGAxFfj1ozWzOYYdC6FQMdP3V2GrO9FMtfY
59D9UC/hzMNoHQOOkuOJa40AV+EN5jq8W1AS+8f3niqaDUcQwbbfM4GzWZyZo96V9lkoul21IFWB
S5ykPb4I35hTu48uYsGa6bciRxEoQk9267GME3eNFfjcuu4uQMD73WrsiSYdC1FzNPjpsHhPFvQx
PcysML4k9baSne7dq9RILCG+wIGYYtyWlK2+kTvyF9CIYx49CPGLCBuQ7Frb4QQElLrl1aBs2+OI
Pz/vrRT0uwsay6rjxv5bXSf8cVSy/fFWXjQdgblVy/bi17hnUq+EP+3Yz8plO8N4N4YBGbyGsRK5
ZOULdRt1ITJ0vJ4gaOlNavUM01jKG4f/mbxXPsT1OHpXsmWgoel68hOE/nGp/YwnawU0YZCW270H
cdOXQPYPEW/UL+OoATAdOx3YEZAwz0y0tkmpKlQ/rTdX1KdTdWrt6qYlnJ4Ptx8BDYdN1vbU8Ux2
YEjlVn14eC2wsCNnV6PCwEMlBHisBtHfmaZYKSrUSX/rIJm6LogMavtfO70Vq3lBje5TViUDQy6Y
RyS2mU2+Z7ol+c4ED5Hnhs1c1GQ2dTOBsP4SBQOidjnKB7+UQHSo3b8q0u/j3kUGnNV3hcF+E/UT
Yf8ZAraANGgsAYUZyc/VSe6pL2AOIt6youY5EjNnmfR01WXgS2xrWzS+ivW1zdRWINldUHGBsfdQ
o4HdOe4hupfIdkD5NxtLMqq43C6Paqx49GUlmfjfSua2FyEzGn5W2yNHnQ1tub6vGXiANDyjIsLt
nTNVOxGy7zWEYwXmfYA0iTghdEQQuPd2UmC4kkt+vGy0fLSiSmRXA8M1XyEIasl7WIQ85ZQiCybT
shnEVAy9BBs6L/TBhJw1pNLqWrQV1ZuERcGo8aX16PIZ4PXdYpjIe9VIlwTYDOWcROodYxxY4XD6
sO5RlRK8TK0J5WmFPaw+MeBxA99fE11iANaMRL+V5hEbgxWhyFKMz2qo4m75JpUcFE5MVFWccPJK
6bMeZ4J++yDjUnlwwO/ffgM+VlfTpDkLMelt2JBJsqlof5KhbESiZ0TVAoyF0cC+8FsrFzy6TU1R
IkHeYi0s1gzebQXDnVpT3isJhmuSSfV2ayU99cCK+U0aQrERhN6xMWRVzY/MGiO6MlB8+oHSNogh
BCVcgjFaLvKP3hceTmKM9WIjSdh3Z/INJJA1/CChpTo42CMUj45pOg14b7RVhpbDDxoB/6dHtvDr
6BL6AYk2HFE+NCELhycypvQYtv7PwvS9RnjqXSJL7ydwyqN8udSQHM2erWWCh2U0FiMrIp8QaKGs
bPkfUQI0Yah0vauYgg6KelpvWhLUmzDe93Hle+AEUeAf8QwjbyPNBNmAg6xx9KZSF9ON8zz7u4x1
+Sl2LDYD33Y+DFrZ1sR6OTp80JMgIgjzDprwwpEggwUT2XiGen23bEov/y8qR/KpmvhazGudZ2V2
u2sT4ouaMDpxw05mOLLxCU+Nnt/FhkNcKXzEUsiKwuQoSSwzCLjnq3pZhTz4s+FPDk6F2AaUq9qe
KJ5CyPLdpSUc9LfhyJaSo7HfTw23jB1YYCWlG+NCLMQftyZYkylINLOrjsIdjuV+5y0QEolabJaq
V4aAzq6Nz2xfIqEbqIZJaon3tZv7u6nqBpG6piQk/vTZhtB5sOQB1+dqCV7t3pIR+ObullGpmHlV
D7UAOPFEKuk97pn5Pjed844cvIC5NgxaTsUwb5tF3tIZ6YYsK1P7iqpzv1BxL6KNWvpjTax3kz0W
cycuq7Ve2Nh1dBqmQA3P36run4yYFHz0Q8p9qdEqLgsry6g25L8cy3qNdzWjvIqMZwyNd658F41O
VlHtRUURcVFtHuSUWakBAjQzSLshGrcOtvh1QV8SnKl4FyUqUmOSHFWPXVrbRxK4wHLa0rYzEhmf
ztaUmLwukkoKXZjLsabsekpHV1X3HHToPGbAG1w8T6B1HM1Rv8NsdIoeTlxASxhgTT7Wr3ZTHWpY
wgc4CDmcc8wpjoAwPsTImtO8QjsNAg9XUUrTnZMaK+BkA+y1BmrEqotpSZgpQ1mt6BPX8sy+SSNg
djTWzIEZBdPqSLS2UmPQjB5YphAuZN2stgYvaDc7eRVEuZn1MblbGrM/WVpnfkHtSRGbsxAvGYdh
T8IdlQlKcaRdHiovYLkVcYeMzwkvI5jAy9JvmASOyVneFCdnC/be4RfCXOjgKHPi0u0C5up3kic3
tvhpJI2jVg8Fx0+uFnP1E8es/EXPuOzKoCf3X5PlZ+/meAmRFecHJnv3H4IOB3fCrfOSrDlKdW8s
I5oXD1Gp23MDqG4W44m3SmqkQtPxUjYeKyXsDdA7LbrKKLRZtMvRpR9qHRkovgbdmrn2C1Rim//b
5rozthvQVZBOgYzO98IWfCmMo5T9POE3uFg3VTvhAcJwdQxoapY3DbofNHWslh+qcKIA1t4zrKFZ
fujR/fbI8Qfr9cR93MclGjwyLj7Ln3SLJkQAyE3AhKbTc3JEsWfsMPCQk1AI4LKSCfHBQHiMTCq5
gCxAjBMW49wfKrHj1GBeED09vfm03HGZT6AuIe+XVnpo5+LUpfTT7clStkS5drIlU6nByHSklvnj
szG2I54zXzyeT6zG2Qca88XuPZFvfgET0oG97KOkArvOxJcEVgb62lZh7kJ4FKt+5AmPRb6gxXQ4
uXD2rTq2Swaxh16mo3LnhZbTGAQWweowikNTskjhWaGqhycboniSTkVhwyHnYtlCm0KYW0p7POOD
tjXQnSyXS1CNOSACZAyRh6l0meAwHrgqTlZmq85h+ni3pxDybhWMv0VQ8tR0+VXEoIN2iCqN0xRL
xmdHn7921NzC03cpmTMw7wIfApOpct6xuWryCH9krcXY+Y+TL0hhJdQtz5aSJS4gBSUuL3b9mShh
FBndZ6LpwXnsotjqYL7FozgyFNmK/7aVHLug+KD20OfadfuZgaL6QM6BoqdQZOEduL77Vd1KbI39
S65qPocYfzAF19lAnd8e6mSQ3KwZlMbYnSnFHTY/nJ3av7Ql/LZu9eD93QnOPM4V2KP0YzsACfZQ
HGpC6N/nZF1W4wT3YHDs6Ia/oXu1U17y36hAGlIVKHnHtoEiAqQz1lTFNW6aRlZLxuNTtB3j/oHd
AUPScSv54uOoaXkC90s7e31fIHoLZ8vWbhKb3tLuRSzmk+cEUUWNOJQBIddsd6dl2oX7oI/MCf0m
VLqGttQydK87XUna4aa/XvR0DPnQ09a7zVzceiOUwsCMnED0q59v5tBB6sh0fPadHK633Fx1IxD0
dcbZ9RxurxYodLs2QlrbsOZ7bheHo/BBibP5OHUBsoAQ5KggvMyq01wViGFSnaKzWA1ell5A0hOQ
tJpChC9gK81oY3CfXd353T8tnPxtprYBgS7M4qXEtL4POctkAx3NjYHaMoE38o3EW6FDkrvnIktJ
N6BLHit/3nTVwyMlEpkDVCPnv7aKsAelqvh6s5bGL7L1ewobldDx9B5FF8t8JS6jC1S5ArFaXFVT
eNDcLUoa22ugNWrP8BgBz74nJFx80iHfaZG2btj8VSKOKv/Ats+hOwEjGoB3BWVs7xxxiyJ8eEpg
KmRYQE6Lyxmjfp9I0MfsVdmZOyG0iwYL5wWIHVPa2bl+MvQo+IPkqJ3qW0FUsnW3tOH0J1JQdhUI
D0csoF1hTcDfrJhN0pyBp0l0N2tA9mpSSQW3YRppuJNomJcxzCbGS4qweTdYRgmYmftqN0HFXRbw
OkhkJN/NiATZAgUQwKBgYqYXHT0sF00S74c8ohd8GMXm/Kid6A1hzGPREDFqmW2g8K6rAHlOjueI
sUkEnkHYNwxYTe7COjETJ+IL+0RYKkt2YhE1DXR+PmGA3EOuDKl8WMR2dQlksO39fWEXd88v1kYd
JwRXr3AyO+gRL5JYUNcKKLCAciu4DZxa1WUfgyzhJbbkapdbqOsxHz4hOevVVy0h2kk5BrvpSsrF
g7Yo7EosfPdGCzD7/iHc12Zb+X0m257cHR7mhUnl9PsJAEzggvzq/47gwuzZIRABhSVzkU+Z9MSz
gCRIB5QAHzGORcvL/anWRpS/YepQY1TFN0sXA01um2pT2sO4K88bANITzvztUTY1AFI35NMYe5lz
LKrUatIDiO4UNMKgMS/38kq5vix8cCq39M8zuX0VKMeMY+kVhuqjdqXh49KWZmIa9JoJFU72c2vA
uY/pB1iuXQmrYMaDP1RuEcJyld77+yY9ewFGJ2D2YtR7NRRYW2dEbU0DSWaWIQqgIeZyRJshuTsD
VYg1tuwn9WIkadGFxrmtMkdNlh0FPi46VxBt9DILGRODgEjQ+Bvg8dhW1oTBx0jvbec0HunGVUEt
y03BcDvTSJ4GZ9Qa4dkBTV/4/AV28DsrDV3lN+QSrDe4JKCdD6HTlkzKnNPkIMou1XL0w0mqopCv
j0EhK9qo0QcYQ4iuMOxW66h11c03NWEgAoV6hlrcarkSr8giQk9wE5UYZnKojC3x8QwlLU5ts27Y
z/5lSvFwLtGxiQfCMFm4gbl4XzV8H9r5DODPT+BUg3KglCW5sTTFg2Nkve5fpZid7Es2ui+yKU8o
h7zS5bzrCIg6MG82geTe5jRoIXI81ThhJSACtaFxGR7zGfhgoEtPWOsv/aBHn9RdgF84TpnFR/qm
JNKKdi4DQN6H0yWblylREa+wEqMgr2ARwF0Mi4kyDbJ5zwwO6Ts1C6hfg5o7NWJ4W0zpS9KuQWBt
5/tAKdOxxzTyAnIq29x4FyemrcxjlkfRTcuyT8PFRkd9dobZ2F3Vkc4D4OV/o0owZ/0hQPX3+s53
glgBjn8TYzSVFnG1yPa9uKgpYUzH2VDxY0vh7F5VOGE1pN5HuB8CmiAqHfGuYyYKBnXQcdSRuJVx
jPB0jC2IK9R7py60yKIw96W3uXqp+cypLP6n5CtDoxhlhdHWte3FK/ASN9gi2URONNFANXG2Cj6p
KMwyVNUpQyGqXfea5zywi1f95snf9330B9o8W9eNzJV4W8HbHY88ec7pscXOrLtjSdr162fkF9uh
WqK/M7ue75ITyJ24znARY1w7gL+Eco+9y+ekt/55X3PZGeNpaK+dSbd7Tb1/YLxR7qWgHSl53pFm
5mEdvZkyO7tGsZw7yaWzlXmunCEy3giQo7wdNKBZJdoW5TrRYTNA9tCldvRUVxRQylVxD/FXs+Tq
2OSMuwvsKaBAReCHvJukDNdQ5z1Vm40JdvQy+Bf81x5va8aIwvBd8eoTOfwuLQRCjQiBoCA73HOS
XbjBEtT/B6HrN2+kmKb8z3ZtIom+XU5tZLskQULty0b2O1bEI0wvSkLL84g7GmQgK6/SLHzu8kfh
m+/Exw+pkWP6chL9LqxCVrnMq+/IL2h9D1sJ/GZwVJZ8/D3JXEQT5pkDq/pb+zV7U01lR4nnYRxy
7hSM1h03fr/6fTpkatym9qsnc4C76wLy0vUqpBp/bpUgGqGkuWfUJQEir/BwJQgh15WpTR0TAdrj
gsGB3vP/py9fFhwy9wOpBOVAYkfWEO4r0EaFfrlDW4X15tX333NBTQy5w9+oNxy+u9nRvlOgE0qH
0eifnVc+HDzce1QR3rdk7zYENzQc6wp+ydodPlABiKVaC2u5a0nQACetJteMNz+z02TefutexRQz
oq4ZhcXiVNpY3kzHurNCwA8RLorlAYZ7hP9jnF54x7M6arqS4f1yDuMOuwG6OkU5MZiotOlio49y
Yg3pT1MzeVPV4WVH5B9EoD3yyZXJgsI98+hZZHzaalNPpFFncvbJWUVzmX7XWHHzB3aVyqwseQpw
6ho8nBi9OKVp7MmKdqNOB/AIExZs8lt3jpOe+8nzzVTg/ArYW/0sCMFQet8iiDgxVLCrVyt3QLys
sszBSDrT1NbHX7OLiFux+9UsBiMKYBLb0+o+QeFXZviaJx2/pD85sXbz6wKNdncfpyi9v8SQN2TP
5HShZUXU+HuZXdzoHU31lVB5R+RSLlWXeJ4V0A3jpBteFXw+BmqnYTtClply2az4iMNLhzZsNFHu
ufqbzofNzr5qmJRqvaFCby62TIk7O5niZlzYAIUA8eeElayv97kz7MkuJQndPso/HOOok8HgZVpL
Sm4ei0qSVJE7hajZsX68UWdD/WoPl1Kf7appuUItYN3Hirouh4ZA6OZcqWk6v19MyTy/1C9UmNDL
bfpNWtj654L1xg7Bo+VJVHdhbWVnZDlPIfi9M80s7ORXxLGacN3mivFiCsWnjNrpTtIHBWZ0FUZi
CQmb8QAZvhkSELSCAu4W/fIiMnmQ5Fg4+e4FZ2fkZBlLSJh7GFmHnIQHJzC6T1xIZ+EQYFwaOtjK
VZljon4ewdx6rBrFvFx7U+UK0m6M7h6mDDSVp5lEw4UOfv3YboRCX0JtW67Tnu0bisGOYtSv+1Qh
bbGq3gSbES6QlUwiYijoTeyIiqt/Nt3XqPHwVCBhxC56oPAX898ziqdjL3Cs/KWXXZWZbUARCDjN
wbubY9onxNZlUBB3RPsE2C3BTzflp+dhw5ec1G+V0P09kH5+yhhnbzpau25Sb0jheL4r4kfByrgM
OXlxPeTvZp+hTqUIqksuVjZbgJq6OJBvNw+ZJLJMJr+oSkj0IInQRUjhwRoD2BJmEu3gJfuUUgpS
WAs/eaKzeBzmHUdd3jJV8wGg4gcCL4YjNLdxLQs46zgOm4dJRmaHjQS+adO/jEeqahBmwxEmkka9
cdDcZwSIsHA2cgFQhctSYUQrWNg6BMKgHJ4Q8oIeb4cIq1U5hWiQs416jWZUg+3GYRxMVaHmk16L
3yDDW56ildyoDnChtCjTdnfcljANfgAs5zCEZpo0hDklyMstMHoRRYT/ekVIv0xGm5dOgAacOqwJ
62zeyRX1JwWvHTQzZx3jtSQjjQbPiI3kHz6Tqcf/qxDJocOo8AzrNnse+MaeSaMVFZHE9nWV+gVG
tm2Pi8p/cIhHr3LpMaSgJz5j44MpRfu7KfHaqSJCS3ys5av5U8VIqRpagY38Wd3xKrpiHNMo4WQC
IralpLjGvsgFwmblyTlLsX4+4ui2ELuqlVmTOPUIX9vxgKeRDOQbpdKgcB0T5zK95bTY+fg1AMsB
jA5zjmOvNuxsorPGopUvfAUI0xDCe0seFdW5Ic0xKfouIIsjC8mqN/zo9vX65BYAAVk/N1N5NuWf
HQ0/OtHflCAY4wKIifSQ0DddBlSomCB0dvxUG8+NkEuml3G/q7ZaAHJdO9xGrQtdsfxXmzT7D4DI
OJSGZ9dD9Q84d85jyVrMFcNLrBk/snGahNwuX2yk0aDA8nQdn8VcGR7laHk3uSpKfXOEz++mcbGY
aQgYCM5y1P1ZnQl09z5FqqTHMKw0xIm+7MPav1fQb7nazfTLqlw5PmBbUPCglHnr5AkNVT/bG082
PQ/qzhADmlHlCuS06kDEBcpxB2Vpeqi1WTApN6jCHmft/W6ZSi15jkw71WGPV5/foImsxotg1jwz
PvfGkknoYBGdKqgmiTVtw8dBnvGlAiWLQwP1q2e8C+DjQn+lo2Al+pFqNzfK+b++wERSnaJ2bNHu
niynSUg07LiOqFJ8JfrmMn/6WqmGdhaLWfD6HhMoXMUeB5Ck+ZrWwCKFSYEG40O1JGJkh0VOjBjo
G81VYmckiWYePTEmCacEzFyNFYGObJfF+fRCdcbwuO2+T3Q+uEgoxr9iuRb5eztEpYBxfnfBgcD2
ibFxTYoKnp6DhJw04436QAf2qs6yLu36hGG0dFe6SzabM9Mfdw7wxrHaYsTIf1s4exYK++LkUb84
CdCnAIzhJyqw3FdUz8JY7fbGnzRQBhCuW6EIFtedhjzpA7/DXNKY+2gYsUfl0AsNQrBtY2CvCuVp
+hXhhD1msDpiab4+LLq3Hx4khm+n82Pnlf/CFiXAItxK95CGNfy/a+dpACKG4D9k0NkeSKQoB7W4
1JRvro33V/kLBjo2j+1DtBjMmcg7/G2jrbHh/zHtKAAkFp8uTwPEuffP2A93dlwT7bD4aoAK2Ttq
MyzabUNvIIOZvKP9YnhPSjmtWZIOQPrCert9sch5E85Qs66XAD0wq29Z4+PJkk6Uq664oB9tzBX9
1SlHvU+yAikEy6FRHc9uMUN6yesGqsGyQsAaVHxQ3MEPll8EA06JQZCN5kPFSdIi7DXLeOJNcvWd
F45Xk0m3NWLjr4Dh80bV/y8w535YKjOZwgvXnGhDKRizA4HlUm2Gi0K/NdkU0CjMFThYDX7v9iIi
1nTjb9H2+1rUD9sQu4NPtM7wTwcK44a965DNp2VEhr0ujBIzCga1gfwFNCBERoeOB9AXDU4Lw4P6
0PQTo7i/2cyop1Wm7as6Z/6NNPk/bMz1nr4DyOJhid2s48qQ2+dSieXzw5zpR9ci5vYx1wG7Hp/F
2Z13HLnmbwKWY1ZKw35R6JCCsjSeygJiaXDZYutIc6ucIKJVxLlaJWYr0JbE7Qg2EHesSK+4wyvE
5JA8hu+Strt8N2Kx91Sle0JvW9GxDyVCdW2ShWkVhABM2hBGIYkVcG4XFVVHjla14sdrATPXUb3A
HeedFdQPRHxSJYOHuhxId//MO83nJqoQCo5qH5m7yt9QXKKW7op/qj0yyXNNkmzUxzvjuW3OQ3oW
26S0DuQbvz7gNRSqMZZG1lVXABjJpLTlVVGUXWxE7DFmh1ZpJaMtzvqZLO7uOfOk0ZRzzmKusSWc
C6ez5UveNF+TsdccusJHoeVOiHUU/M83ZtkiKwOX9kW9+VJOyyeL6Qzi+vVtBEvVufmAyzavRXxv
zy7NoSkMqleIpU65eRHIMWQf293TuCOWL2as6T7W1jwJVXN33DBOvmXHw0GgWizoYHLZ2oVs6aX3
O7iJDiArDqeZY38/tbvqSOFQHajLkPvMb+QnlqYHpHxflvNq3T8uO7QaxTQ2Opi0oiHKlbLo+aPO
yYlnRXa5TEjo0VtFl8x3CgD/Z9Nstz2xSb8VAgPMYvMhLBjth4qPo6Z9QCeTS0GTcXDmWIHgKet6
8n64m4wPQQ2Uu076lQrWvHDFZm43RKgg5JojIFjubEhR2OFOq/6xLyBZyIngO6budrDY9JJe2T6T
P59VtPIx7YdrsK15kX+YXHBDS6befRcw90N7vv0U518jHhK+vtglcWKPnPE16etX2XmuJwVlJsAQ
iwLggIl9Q3Cxrf6QOpjed2N+ESJU1Bg+sNYVacZbe+DdlT3lxxmwOo6bN/EsZmFBqMr9i/ZdcvaD
7EszsCm2AavLQtRt04TaruCp1Vu7Fg0zkvskijzfWj0jBuqmQyZKpIOFwnRe0A0RiIO20Uf/mH5j
s8Y8rKAReKBP1nTjlX5ytm1DUhio1Pmo5sfnqwz2WVchc1/hhhpS+UhFCRweznA+cMaBjIIhT6Fk
McnC52e3jE+7o5XOPD4R+Y9z2F36E7SGoH4cR6zff+BqNM6OtH5sTIjRJeKtUDEoOhr5VHhROqJI
YrSLabihgqdoQ4gYuUAYeaWAmwU5o9+rMpehxNTostBiP2fvtl+oWjGeRDlWFUviFsu9CvjvC5mx
PGg8bw4lSmzudRCx+D29ShRVrS7ynxWa5zda/efQbU2PM45jU5epGY99uvy5r5kCjyYfVRKcWil2
4DXa6akJPFlWtQM3rcOPhz2JnjI4vsnrwKJ+78wh9zkTGcQUnEZtN4LfRcW/B5Z5MPIrTZGDpoRA
32NoIcbLqUvo0yVHeuRrPLvOE6ZF33Gm/K1wWc/99SS0beD5Sro4ET60t7F/PAqQpln0fbBkcT65
TXzcQTPnY9f0oyYdwdcdHW6meVPXUZ2Q6GLgZAV5HU8E+2x3ess6fIVnPqjPveuzkWMjA0WegvjJ
825nhuPh6i3soctSrVli4msi8JD5wYymxjuUIR+Pl+9UxYDMRTqWxWI9qkQcsCNSi8WKW8A16zWF
LZ7LiuvwEmypYwnDJ15dbTxtjqcb24ybnHTHduyN7a/P0emt4GH8Dpz3N4gKuM6IejF3X0CmHYjZ
s6pWC+QJDkxPaJ+p7Toz1qQ3K8OM+FUKPg4aa7V5RhG3X1iuHLSkUsNuu/0ooco2+MRs3/G8zUlO
I70mexalMY9qiZpJDMc9AyU+uKMewg+BnAoh70kR+gGClsz0GXBXmoAEqyRjx8UQ0lqRPMn+JPd9
2uC+uRbZd1xzYJvFSkuPRTaqxyrV03amqvVu/okdw6Ile9tqNmKMae4g8x6/MhMtkb5j5VSBfiUb
kWxbm4xE5OD0AxLV2gaAizoyjeJSM5ksbT7cYRjzrIHy04CUsJ9/3ri64zy+DHXmUzXdPoeduD7u
DXk4WkWJknLhDAWZhFsw/NzBQxEDh5si69HzRanobc7w+nxb6dRo2FYL0R1NXl/sMTDfMT+HwgK/
XJDI0r0WjhYp/vOCM23bfOK8zEWlxmuldE2c6KwlUav3ULmtkpRR+L43R+PeSLcq5h5d8XS96Yuj
zYxMVNnxOXyCtNyZEPaL+WLzhpBvFf6O8vVsVY8/JbnlKa6YpUEyI+qNtYRRONkCGtxYwfHy4dDL
RiP/F/2Mx7nenoeSlX98eduOuI1GwpIk1+ztGmIlM9lK7DLf4tmOSdPIz0K0efbfNul2XHrg/BxY
Zt97uKa8hxW0Gquj4sNdVOBRJ1Q64s0LwumbLM77IXPa3CKYH/XKVljkvZYYI/FjQI26AMl2pU8G
irq65PEgHCkcBmF6wYQ2UUGkILNz5jiTY3loOaBDcz0ToqxR3wbf4kBOLJtimZ0jH7dOf4H57Nus
Y4eVhC1YCSoAaIip8QoGoh3Z2Ah0bL9blo16+tlIJvzWzp4pMzjdqFFuOn595mWfSBnmp3zviDmn
IfPt1/7zUQc0T8AvEfDsnUIk2lOCD8QNVQ2mJAcK3UoRARa0W2yLM/sVhBFPEr4Cn2TmzdU1xbtb
OHx/mKCGHvHwWLQG9Rp6DaMGilDGaA2wWtM2JTwjRg0xcKgqvkjXVoatwBYWzypXXKYBW4bdmohP
r/SLJe1tM3R2lCEJuZEduTqOEmuSxfuHfV+h2qVCZG2evdgq1dCZwjhNjn+FcuFUScQE4Ag3eULo
pv8jQFlyMqnYYexUp6DOhLx9T9nz9OqHHEoMTXW2J5VETS1m9oWPJyAvWiEIKFkJqxNjWcoWD7Ht
PRoVZfM4kLjA76MEPKe9n2h9I8cZBcdBfLxKJgl77voHAV+JiDTdxW5uY42/bh8W7PLA0y9k94yh
/YzvTMKrf2k+TCnw4ZCyVTQ9cOosPaoEmmmSfXxLQ3bmyfk2tdCE/qwZ9RAtM9afPyxEyQMs0ya3
Rck11hbqHVSkkMY9kaeTVzxktVisUo9FBdM8u+v4zmfFjrWTZRby82hY3BruGkD+7HmgkSBoDyIP
ToFXA94Yv5A24NdXANxtH0wVvlDk/yQMVgBVyGfdMIPOEVNqC1rLIwJNkg/n/6SD24fysEn7Lgau
iVTR7GRiQV57SPb+m6Ygyc+ipQbfJtrqG7tMSPXt87gURjmufMN9rhcsQzFW/ypFvN/l/lXeQLuE
TYzW9QQRFYARrZaeHou6VhvEavpKeeJFKQ2j0HoL7/sVGmBs4G2Kx3t6pMA59ZlsQKuSQb0nt5S4
6m0ZMgDKNYV4UEogYnoKeiBgzppw2cH0ozILUskHylAEN59UAGi4od5QHrB1wPl9zjocOx3rRBEf
y/JqHxbeTXUsSTaj52HBo0xy8/jGrbA098nSvj1T3dabMv3ULAV2nGhSfBlRs2Lc9H0qmf/EPeEZ
+tHm6jdJ8Zbm4rKZXbqdhzNz7FRingt5XMhs36zI3B5j1MdAsCRc8nEb97cUe2LF9miOfG6zfeqL
MF35ww1K7fUarDST6y4JruI+62e7Y940G3uHZcSEpRBmCa11Wsb8GdIsODqpDzb/tp31qPC4LzKO
RlKhjZtQyHuVzvqcdyKNY8SnwEUiZN+5MDUSKJOoV7MYGGeETOrBxf/u24urFJOj4bY/1QnAkx3E
aF9jpTlu/8YdjxiH5JVCcrEBINhxHurMLR1XmOYreiJLBpcSkWH7kH7I9iIg6xwOP9O3+xk9qfpi
D3FJVZ8m85dmMG5OPJTu7Wiiu7kqrQCe8UsJM5XNDGB+tBOP+xyrkAeNz6a817h85ZUjOwqpcTJQ
+PSNEYzPfcBWTfQ+R9PbL1D6fCYehKBfxo3xt6qiN80n5Auj34Bmd4h3303THoh6letjjnt8+XED
PukgO8hQj8vCGp73MvvlA8sdTok8DKyA0ySHD4vInUUbkKgWyxKIq1zbKaiadAbl2uhmcwXUxftV
xgXi5W+L8Dx9adAMHOmqXEcT+NNNV0bqHcycZ3276B+hSVLZRVEO6CjJv373t7hI78UbTTJFsjHh
QPGu5iM9+JD/84+2gFDqWGzO3JTLOngF/pjaJAnzyNxWZ/IqWkWnW/9QZTQDE+GC6e6NgLY541w7
nbAKZ3tKpekBXcCBmRTFmlkWJ9MirEl5TKUmyPVBmdd/smILdCK6YKQApdeXus7Z5P0Cub9eZYsV
AZToBDx7D4xQMvk7Z5hgtC5OP3D9tX4uGiOpl05U3EmfM8II81qH+mpu4cjlnpaR8EG9xJoYMpl2
vSZVz6erdWPHkVKlAZz9p+nrGTun2xUlzgg8/5NsI0AlHNX3jD+L8Pw77pm/klSSiOUr6qP4A/1R
/aYHniJERsnm8G3Uz4w4TYS3LIrN0no4JxdZZHr6CQeQuhhws7fwbQVchqE4irAO3psdTAuuUPOB
3R3nJ2K/BGJNxkBVIgxaxzYcV4gY6dlGnF0lm9J0u9uTj9pAH+5kcLVj+sIlm+3Rw3GFjHEJBiDX
nRjOMY9CS1+m2uTSFgvlM6XJSv9CAGSHR6xNtqAGvZ5IANmp3X89qfz7DzVlzGsOIsEOd///nM0b
Bsj8m6+cpnJ+5zIoHhUFITg5tvfYlnhB/hlAsdTVnlASKS7uEZC2GLVWXq2kqyOsEK6RyZ1LWZ3y
pDAQEshQAE7U4CJVVRiFDWorIS68gFF2HHmxIKrw4VA9D/Weye2Dc4dc11yX+eLxl54dOcc0dZvy
Ekv5NGaIEuGFTh2qDCa2SxgSqNcWNGTd8SmtK0fMuPT69HOQfZ0IssSH33Vs3sFC8SDobDj5tdm3
y9Y7/ViJfgNTVJbOkaLk1IrFWnBWyiFM2n+cLQefcsiL7xPM6M/QUDVKRVbXjYvLzwD4LqJIjdrU
YS7s4Hdr0oali9zJI85f9/WE/nD+CwJYJ5eoei+Qs7avCp4Rn+VVPiqO4DneUvg6GxhRginZl8NV
SzHhF4i8fkpktOhOUPp6CMA9gwNUCENtqbQsuEd9rWVle8OVglDmAbSY7/KVW3SGmMs0Ycc8oSJH
FbLnLX6IkXbkpViJ5prSAlqoFATSFqGdrP2Uo2TBkuENFc/05veHJXMVBCqDd7AE0wQD/KdldUnp
qReaGu4F10hxYV38S09jL4pwqjL3ZdGtFPuKHTyOUSH+4pZThEEGdH6IMg27prRINAfKDpBbd0Oa
F3Y26Y1Es8gCKwU697YwDjT2hlLlwigsh/Q5MKOe0nlA6WbiPxcjhY45ttnyVZfskO/qtfaVIuX5
lEa5cDqxpRopfHXmtcdWlKVpNJ0mECXqv6I7jqbAn4mBAjeV7Y2i/29C0W8RX5a2lzHsP0miXfUg
U32Sg+yLCJ7OlQXIMOUY9fa1fOsEm7jTS5YyneibbGFr5QwVcfhC9i+tnCaqvxuv+/6zv6mQTjJG
IZIaINPB02sPHBrTATVxiGoze8typS4HFQTJm4g8ow766eYEf8ZsuBw8cKA7srxkjmY+SBVQiNdc
xVTxvjMw7QIuDkRcrT7PSpnWJl+IPh4GrXXbk+aZZ/eyohN9ordS4Btyv4UnGqtSJuAc24Gb/gnz
T7ktmruwjJybQxurbJjwTKVWM6Ylp/qr/mKhoH4dCvjotcAP7INkE22NC5FXnEju6GDJZINk6QNO
OSJaDicFX4uZsAv8Vn4L9ZUEvhEuZ1380F/kqtBg+dnBCjPgxdiw+/sC+4+tJi+NhvZLxOgCga7g
I/j3+1DvyZ3/FBQG5kItb2/qTDNL4s6jTaKG2FwLeAZJWE6SRV82rtgN28g53bDGCpLGEvbhMwTf
DUAFuPnHxxT5iC7xfUhgWvBAHoA1MsQ4c2DuULlSzdzQ9LN+vFH5on+w3lTZog8CGCcEyOR8x8Gb
0ds6odMZafUlFPFxXbY0wt1UWTJHwmQioCC1GUjwFJSaC0TNgAWIBUdo85ukuIl3tlV453BI7+fX
rgm9CzuU/22AocbW5bNuEEkZbNWml/+JOCKgptVdglbJoRxXLbWjRa1XFCvY2+vC9h2BVmeIwyLZ
ry+v9YDmUqsYcHt1FRlfHE3HGLtEU2RbVOtwo0GdiBeRHa5LIpm3Jv3RlfnToF9fVl8ud6Gzre91
567085FuW1m6FsQ2hBCstNxq/M2dA4WPPYBA4RMBIW/Q6XpccdAzWAjjnWLj5lujjAx5W0RRwz9I
MoTlSspsR/E6DhCHcfMnAoC91U4bLF9S0BvqDbjUfIwFFiL+R7ZLQ7cQWXarC5L2Nmy+AxGgy9Z3
PB5BHlf/dix8TLSeOhtgB9zBOzuyi9SNIl5raKwJZC6wvlZQu3d3WF7kX/++zrIdlucx3hNcpHlw
q4mtyBv8U25gf1UR/BL3Ipy2wKMslT5s+bH5Ks/oOhiyblyfrSs8Tux7Hkr3ARTy3ol1TfyME7hp
bfI8f2CN5ZybAnmU5wepkfKv239SClL71n4GwXeNNHODbIMcPSzP9KKejK4flwKqp9xdyXESeNaN
2JRMXX9bicZlxT71KOkeufIY19YLf+IBXYqQgo3oDBmRbSEQhh3+JxEk6+mJ6usfTKNkxcjnDoHa
vaOqU1xXWo5mkPvPFR40ZkEWw+JCPFMxixP+8qPrlGSEb1yXXM9r/QqNJ5TZt25omEVFpQHNcKSx
Q8d9EnKAwFT7yiv6Z2U79sT1ulp27A/5As5ezOe66M5m9tAnD8xEyK2BvjBZLvq66Up7DChTLENS
FOWY3b+YkFz9quRVegjYuwRuLa2FgC4s3vH3UUKYa6DhTTj+84bPHvXNgiS7QDpZNqb4McNIZ3ok
PWS81mL4LAJaJnRebGTsy6G61l7DH4sLTF0ADZ9khCg99BCLDHCVINkfC1VPBXP0DdSKr8Nr9J1D
1xydhR5ilkyvs1gxgvBGBQAYuxCfbRgHO5h/V7JtlHZ33RpNEApmMV4yaRIoN8IVwFxCuxmMGY7C
eJCeWsimxlw6qKGZm8IOSe63K2coRjy5ufUq/x+/XFVwkf7LiPJmR+sKqQPj/nfy389FTqRcdpqA
uiOLKhJq0R1TgKW4iqac+Exxecd8B7GncmEdMz/Ns/t6DafJRtb3v5qAY8pDccYLPdqtfO772oPw
CFTNdrSQ1EqBdjve80Ya9ktxqK2RnT76eAyBYmq0rE+M4/vP2BbiWPohzQ8bZCDdof29XN8M99ov
IsTVGd3tomQVPCa8N9C/hRt5kg14wsr7xSCeC+xizbek7NYC+JqdStOfJw3CY7JGcLltcxi4kHjb
+HHBxlCFDydG1UcgZag37OdzyxqhT7MF8uZSmG7jiCRl97uM6J2zJE4LD29vSbvdnVU0IoxKFxap
OThLcfNljMtw4nZdRAAbVYbLbGNw/o/G3/QX0/edcIHJDI53bLRclpc69booTfjU/AyShxgfWTjF
dWY/2fARDcmubfQlcdnT/5nmrkUnLv1AzI+0G/mbpp432GxkAK2CjqLZy7QQKXpUfnLOzz6z6SdP
kqcxnPsvNDxvSHwNR2jWkSkODXJGJMFR5TfZtOxDeHHNrE8sPMtr475l+nMA/A2pprJa547MsMnZ
TJTEpxSyJOOMI/PdeP3DbZkoNJ7NJpcXFB/yGUkObD/0MPbxB1fnBTIOhYSNunQiPWRjqWqqSwwr
iIw0E2gxFVbIQSZnrabbksvB02rOHucH8bwgoYVcEUR3ap2Ip9c3YFK1NhKmgpwtVUJdNvYPqzHj
DEi0k3HmdNE0wBAsHRsWWR+kH1Ntlt69/97xZxHffQ4TpNa36wtWWqWqi/Z2FPNOKyEVC1zQ6htc
I/6xKAzPrsw++9Pk+gVavPWI+gny7a3KaL+3Dfw6mJl1TbbmW4V3gBJJLxKdNp9rJ5OMNhasEc2P
HocpFWTN5IsY/h+3LKIYMYwfOz6UQA+GRo+I8rZNQ0szdCo/atx48pYWfgz6wNjYePt7+I39MPte
a7BjjF5NVmnmFdk6BfCLp42T1pNHGBEJ6oX4gPmusg0FgTwuzxwuAURE0aV4qlw5wOBZYef5b13i
ZzQSWrlMClGqphwe3JurbLCwB2yyhVSvE+7i/04FzcpkzeX7SrKLj7ouPeLLnfiEGbH+sRV99Q6K
laV1dGpGo9ejCo1oiW3ZZSY2V97845BTEDSSoFsshuVzbBnaXxLvS0BZ4mTpKwoDczo5C3LfFViE
ZgUlVIC2UQ3CAlxaCczEhQOWmBhjWD96RReqmHaOz4cMyBMzvN3DgIpgNoZUYGdkt+pb8XbWE9dq
5lc6ENPxSFK0f7Hu2EmsWhCFuay3VsGwyBWt9aQ2+iW/7Wbb7zNo+O5EAKKRgGTKiHVfK4I9z4Zw
fiLGRjCnq3LQpIFBBiP4eTjdPn5ljXvY8RSmdXuoeA8L88Bo63SphIGDuUwdl9VIxFkhE4w4PCcv
nJ3SSPuiPOpSfOXQ501jAOpdyJ3Ur8NVugyiAlPbOiU+T+dVGqRt56M+e9p/ZAoD1Uh4WVYIskTO
o7W2Ftqu/g0TTa6GZYF+Y1uFVgp2AQtK9xwkq34Xp0Et20oKR2KlQHohgMuysrBc1ViebWRZU86e
7NQjrYFi2H05WMvngE0qzftG0hnYL+ddIoKKS7fKEkO8l1T5dgQnOV+IoYO818nk478opWlOHipK
6TdcJegG+RVUMmhEEsh5RMhgm1UXPSMKB01k1v+T2MJIABhZsnCBy603V0cU7MpmNZ4qFSo8VrS1
ng7u7q+6Lzr/fOBx8ViTqU97Z/7a+e/tPg9ZPxyfDJ+wOv+a7f9N/i7W3OvDywMgE4+mcUlU7fBB
RsNtK2Zb8DjLSTTalA8iB6SDdO5whFmb9DlYOP9rVpADOLDHt5dgKT9I6qrGw6PQ5C81yoqx5uG6
QafH1HJcGcqfSdlpmnUKtsfUwPb+o/JZ9aaIZc0Tb4WfLBBe77YzPeV3w+Pp4O6Mj50ZfPZ8LL+M
Rhq336ZDs65Vcb53wLOyJrfvRK/NwjK3T6TTRwKKOmpDEfNGV0W0q7IpMURYxUAWWTPUkeoscVDt
i+f/1N9g9YbcqmYOGIXjs7Af0r/rVtDDZLh2yxmCAd3saPvPa2KVtC+zI8kRsIbjIFdFR4Ia632/
lVbQ5BtjyR7oJ2YuGnI9mXw7XIDgNLbcdJSYR9k0YXbE9I9lUvCgZwhmOgT65ex3C6ZL3GPbsRBJ
KENAdjyHC7eA4EWMuQ0x/zZ9iI4fy+S+pP6SRfuv59sI8abgqeOFqg2tgLYXeNfLva8ekx2dlqKi
m7JToYuSt0EU4uLGCbWCq6HdYYCDEwRB+qtwWlD4U/cpOFgs1bs9xszth4wuZ6m4x9f+gJSPX3w1
lrcD0W2YC/9Jtcr4RCoQjzhPSVhm1QvG/CYf9SLsgKcc9LdLOz2vyIQo6ogK5RLCTt5lZ/6FLZQu
tr8Lr7ITggiBpyKtaKn65zrLMnpNbFOjTSlfMjfAIq6g1curvE6Sb2/PNip0/Df95RAD7bCCnbbp
VfUy5nXDwhCKK3skJGydSnw3nzsuBENIJiMEvdeqEmFnoq2jDWhwMHqiCX+OShRZS/mVFTv9bnBO
Q9EQ99OYftY37ePZGA1cNlzqAcPMnq7tPn+jwJwgpQcwolBu7utX54Fpbe64RYHwbTzSq6hNQlou
9KZ48clytrYvGyldXmISzS24/PVaCTTtDPFM/q8LB2gbqrvaUYC6+MFreebBW5+B7ss1FlvQ72rK
d+reI3XsNChz4SZv1PINur77ojqj8jGyxZXdOORfgyo+0H2ReWydPOqZ8YKNMzKTzhewPu+Udg5U
luIayxnlbWnP8d9aD2L/KN2D1mepfoo0DFbEBUvN1UCB9PbMdMItWumZo68yqpr4nC3ZLiUzQQ3A
GXIOd5KWZh7fEQv6IxtjFpaNf/PNZqkrUIBjWbBeECTyggs44+trWqTePf28O/FO7IpGCfFpJAnH
vVBOSocTsbgRJeKWc9ePCoEgRLUHJSIEJBxzNq2qrGFWlFtong2hpT4s2IMTL1elq1XCKtsbuviN
ZkKlu5qGP8mB21pYzSe8UWWA0IaaQukOfCH2gvsa/gFCe+R+FP5Xe1Qtm+zQogcgk462JyAaCoiH
jJBLw47vd3V5pSi+XrlNUsn8NVvCt8tqZa4yHPkZwF1rdwh5AZ035vF73pD23WLNZF67iesX80of
9XJRa9HABi3XeEmEMwFoa1TV7j7Tc6R1vCRUCFTJcP6S93zuZ3qW8QMstwI1r8W8qa/WjxplKqGe
jlIQXL3RZBdo58DQ1xx0DxFl3ujMc37Q9VBFHZ0L7hMD1LhqMrPLkdTEaQDz62KSavY7cSIrdJWo
nTLQjlTMAMJWlUIGBWAqk/Ja3Ab89f4YZwp4KQ+U219rsEJ77OYOeqoRaKh4ApgWVuMLYDmQ5lzH
udg6DtgKl5p/rrQU3tcd/C5XRdBaDx4hi1TmFqu1JnHgW/ND+u8ciwohi7/uHVShDhpkKue+5ouW
GzIPtT8xRZVhPynVN8kXE+Y2QhaA5Y7yxHuKVpQ/JS4Rgxl8mJWM2CTRrmhP+F7KFsLofLM5rcfh
ctcTM4x3zaat9FLxUFcID1MyLOPlznzfKgAvkcm1GsaE0adOFM/0+fD6J8qZ5xTCe80/DU07VGB4
ajQCPYks+kRAE4dtJ+qWxiICBeK35XmeEu4hVNeGSdqX3DNi2v9JBBivBdYBq2Wn16tNeH3kA9L1
xnJ4uH9zJEI0Qvcg9tSu+TZhutYisSfMPqo3o6O0BYUXbtrObPaR605YlQTQISUlRz8tYeUo026D
kIW8ZLQ2ahOkNJ7X81Nd4dOV5id2j9DapTKkl+tEEIL4ZblTl5SCiPSHRrlwCAROB4+7U+57iMyW
yzLNhaaEPE3vIQQc3kMnEyPMbrsKpFOu4U0kuSCzjBBb5fiRQkduyAlZOgz4F5MWxUfuDnkjqXaQ
g+cohRLZXss+po1x1+5RnANeHpQT6P3+66T3Ovt5enj2VYEXgqWky2XbYUqZ/3w/iUqNJAw2stlc
Nz2Yb9rVjMv5CrUFIxEeWeYH7LS9Y8AGtrz3kwkkezNY01tzkql1ZS24l0GfHc2xkKYTvmg5C61+
DsWpIiiD0/kMMvt5/MnQKDhhsVbK8OwIs5mXx14CERrzdsDgTjmAN0DGd/lICVA/a5236P3t7+q8
NKiloIDL1DBmXAbdSIv9WZ+b93e9Cpf13HocXihyr3371rt26kaib6mK0+vMZOkEGH2UEmITNRJF
f+HyAXMGXktD8Y5hivOboOv9Q1OPPnIspsTS7zaMlOiM/dWpZramQHO6+o+1O2gwQoXxqEoGYuWZ
AXUUkdxKa/Dumon3rn7OISxR2kshCSQclQAfQTCqgT8xPWY10R74iTat0ALKvUdQaDZ7aGP6yukj
AOyjITsMlNbNUIu6Cq9r2JrYwrMymX+dcThPsBoUeo0tk/YXwGIwvdRKtcLjzTiWuycWLrqv92U1
q3tmKpMalkS1WvKuaatellRV2GQPSjKntkeMZFUzvwby8KTMzl4xsl8HA6kPncQgJTgABb4XAQWq
cVNT/JUJhodJsjZnjgnn//LQPX+idxU26f8Jg+jX9KGBhNQLLK6Sam/vmi9e/2Adp52/n/Vi+stz
ALv8mgTIZlbDQcBAkktNOcg4J2FJg9SWV3Jg+IMSBY0IR3CUfRbBiKbG+tHc02MWvT/3Jd3C49Ld
C4/oiYJ+N3/tpQ2D0HaoQY/vPiT1DdZtnMfPPF9Ezd7r5iuyP2yOhfHYpcpevPEEj7/Xbl7yVUtY
yTQA5GRVsDUD3P9rmHQupAJLfJJi8IgMAPcTpFa/Pj8/4A2TSaBv6jZaBAXrhub1j//gOAv4GR4m
MhtlIFjKWAIugJ1xzkKzBdaOJkbMD29qcEFSQA5x6mz35sllhFwfmOdlX0cXASUoKZjp6Lj9QnYw
3a8LbY2ydZGPZ5C91EmvrrtVgOjUGk819YQdMwrQVdUDl27+5t5STB7AQYaJXtg7Gq8RUf4KcBLt
iwlMwaJrksLluYThn+fyLwX/vxvb2WE70M0fWhnliDLqMGQC/XDTFl7qiBsSU6KgRZBEt3cozA2E
keU06t64W2v7WYa9KIV6qEyX/0/1g9OMOOFd/Wq+p8O9UFG2drr+/2OfQuVt/HOVR/Vp0goYbc8M
ohCMnwZMq1748YiTdwWAhvp3qLjdyoST4nqZIPvqz0N7YQmKqXoNq6k6rZG3XWo4Hw83DBvansDY
50vvaCEhcoIACY0ZDgAGKR/bv5q9snJRGdW3z2LHaFNsnPjg46f0S1I+qd0bEYJEBX5ruDzl0tpk
cJFH3fUUkdnhjzaJ4oCJ0mqDOZn/N9Ur94Xr8YByH/rrk03dMy6g7HUDsABMgYzOuXSN1Xund6Xn
lYt76Czvb22oIXXnkpkWnrJNoAEtYTqEVBLHv6w0zaplofE7OcYtdz+lcr1e4kB+HXPp9ZI+FD/y
+x5VvH25u4iNWNtHx6HR3oYF6PNuSqqV+ZjEagwRGBLXnDHf53umGhPzTxlniKTqeV8b4B9l+q+L
5K8oW1++IRlsT3Q8FntvA0qnN1oC5Iw3P5sEMYcSr43sghanPiIgO/rJR32cP+gJo9cYdCGHwhbT
pNHTA4sHaajSWjop3ZDAt7wbuPWIBk/1IVONztTt1gco7suTyLcZXut9PWSlwLKp0vSPU6fEnQad
+/i4lT94Hs+lieJ+vKUzatO/AcY6sM/LcnEH7KgNbV+JqY4cGniSimAMXN0osAculJ/wfrinHqGc
Duzt5P/waEwxfV1NkiBTcWzIbOCAnU73vyvrkF5vTIS6935RkRu/gcnVJmiRoZdC7evq1kcq7Q5X
bodIckYCFZEr3jClO9xPgIkjfkbJ2PEylQde8P986xtROzyjBI0jsNOtgsU+Z7gK7ejPg4OHt/z1
lGD5GssyMdNy+MlPK4QZMMPDivAc+7h7MAwDz58pLyWWGIn3DSQ173Luah1FMx3poBPws+hj9aOQ
V6gxsYkIXbrB8ZvLEU+vmXEIURDurG12ukVWtwjZi7CRNFGNO9pd2MZTjb/79SsgqF0vHkJbJIpu
go3OwvLb0t6iJba1ceQ5wsui0d1iEOMwage/eqiWHHykBSrNRIAGxGZPs4ZFTY5ElPJJGrLrq5Bn
/JHkaboMvLURdzNBG4UVe2EPvFrZQQ1iK1cR+SWRD+8Bzims2syzaXDOOSgTI/X2V7CxvTiegisM
AcHlAcxEolNvqmGPfMgFlgnx6kZregA06Y/ahRBodwwXQdgJTBsksvI1qD45YwQ96dzXgDj33dzH
GF3sXpZewFePNG8AldJVi859U/SKeZ4N/svOR6si/QE9qDuut7eF0/mhIqDCbBrJl4W96ScojgMn
/afH2m3+PZiMSwLPm//p2XW94L1og5dxPn6ZoHBq5coEFagsnyeB3rG1ErdPR1Cwk1+MqZsKi1Lc
Sgq9XrHUzk2b4wt4fj8Ch4zM7RZWOG3RnRkQ6cXvboQctg6NnE4V6y9k7ro5C5Nb4/uws+SP3FG6
yKVfOCaoab1sHLMBFcFrAQ2RRCWJomguarJfi+ACIKhX41F+jgHEtDqlqoujFw+ix+irxiS4xMaI
6o6i5kb1XAIMYwSocXWex1D7ZHfqMKjzbLLsA2UwRnoNDHLVVsPqXD7JuTrD90y7bmCYF6mACSJL
8hrNg7NKrIwsRyCbruVhF5g1I6a89mEjXR519k/+6xJ8aQ/YglcVV1mDM+ZAkFpMjm9HEfPvwzq5
MKnoqD9r2aE/n36t3mkPXYkCwXL4JZX/S+QnaI86KMQmfsB7q1oKE1ry0E9Tm3q9XYqTl6j1oCVq
HuEin5pHTK3Kzo+21CQaPGMPctN6aU9OoSJUgEpE7lp4IPzYDzLuKuzV+12u+gTpOu0KWDicKNUR
K7aKwpm+xm97OxH8sfJVsuJO/UhuiMC63rdgARV5xGyl0KTrd3VAAUQB5HL/270diV7Aujs+4afB
izjvx7KY8moqoxpWIJvCUf+tO4vjUzGLY58yXYJ1mLX9mxrIQz4Y4ZwqvMxtcC/TuDCw0ku0Cc3Z
6iPEdzwMTGs3xmIwautD1QYoTi3Y0Y/18OXwGXtpve+qRjXk1SL/LWWiFI4kBQqJ8OvMwzaXf9hP
R3B1Wan0TMiPGbTr8BQjGMlXIonzdCv9qWdFpJIPiRcOX9nxCp63oqvuYASi+fuwzRq5+NJkTqul
5TEoLl91MPXLbxspWu90VLj8tJuIt4A+bA+hr6/k1qKIoA0B5gOBClrU9nfG8laHi1dVRPAzRW0B
bhR9tZFFKVYu1vX+x2LV25Sj36M6HYJNTPhbd99GiaNwR5hZgBgsYU2Zf/06P+IAp6eLMLCuNZbg
OMEonXgQt+wmgN9WMXrQ/KLpqkynQrSi1WB355kzVg68Q2lc8tiDAyQF+HCalLwYxddZt64yG9u9
Ip0Gh6l/Czga75hqF57oSwFYjza+H++LpDyuDQMo0lq9J1DDlv+tkle7ypJwQ7BYn686ZPU6QgAO
xMdjTr2bX2eeqcygdYnuuzLyBGzUsAXvQlNM4nsg3xY8ObCkcuO/3hCwuteXJplHqaeipaX/7rYD
+wMzZaTpV0fR6JNghMCFd+XCL6QfjZJFGzt8pPMZTPTBKvpXyBfZSueu9luVRNRbMzPiihASPIdm
rAI444jrikkoPwNJRq4D+JCY4NF6QRm/zjcfeY3+yWrhYVkXCP3q0C0T3F+DIj+OFArz7TbRddTu
DpStECZm1j2kRjKGxd2+Mahblr+h7QAtMuqAZ7TFTVkfCR0WX+aORIUv2MJNTgT/P1MNiEJowZ0B
9Blvw7Gp6cxJdwHBvwfJ0b3lhCA5GFwQcKeEU71Eqh1amFys1kDB7BOWVHQpKyv2OdlwEwVjB/RS
JG+ZhJZBXY+MAuwIfv8jTSx3vB0WjHDQN8221iEBCqfSEFnbyNXlmL7cPu/EQiocd2F1MoOG7be4
qXb/XIPaltNxEHbmHegxK6uyauJE0gtFPDFIHEwf2lUaf4im4YDLtLVY5U2HkQOyEwKmXchTaLlk
615Ch5+WZi8DFT+8Tb2q7BgkzsDN2Ss5XyYVLK7LTVm4K4hQR9FXj8blj7OnoRGVDhSt4CfBtnDH
rbialI2BsNmv8EcMuGXZbbfV5U8hWWSp8+NxmkPbqt2czXmLtsX2ElJ8972o+IVbdnJwsrrdcMJq
eGvMN02YciFilJ/aZ6V/pBov9EpEC0DCsjySSY3ocw0rzSZgWkkKJjgP5XERlLF3TP2Tg9QQERuT
7VeifJZwV7mhidgiKo+5tHUrA9+RgnuzNSJF/OMktXyxT7oJaZS9otzWTQ50+qdYCmcO2xg3MluO
RL32LDEUfgLUU0b+sLFCNNXeGnLCDEH460011qbDSxz2lvo7dkuKMRshHsQYL+8z0orjhB6GSULj
ByqdnNN7k6CEl8O4/vXHNec/UezPNfP/uEsapfPO1i9YKsIF3pcNLeLoKvzg247Eqp1NybplI1oK
qvFOGeJVohRFccbZ7qp7fds/mZ5ao5Nh/eYk5A+ZSbaTH8EXvAHJjn2Qtg5QKFPGnaEOdazOS2rB
zkl4VelCJMzlqKpL75tS+wj19dwU98invWYHLnf4bTM45K7A7xNiwdrSvpoGBcUByd575pSY68Rs
2cvt/uWmQ+e2oN1bADLnjg08IgZ7hQEYBz6Ov9kMjgZcdYSRwWSlcZHIGpzWo0h/j4PlR4rpsJh/
9J3EMgEVUDXIYL9h2SVRPFxX2z/yivRP7yKAUx2zlXPAMJFJFGTcS2m78lL0mIt0BxIH9SySp5hg
KVw/mbZWhdum0fyS3nTx215MQP4eKf1aE34RD1R/K2DtAyoeSaD7/kNEqLsdSQBtFLNcYovYr5DD
X4dTqkroF2+A6aOZwcfFgw3UgYBRJIuV1idLoklduBhfP/EGEb+gpl1PqJZZms31bNoaHnqrCsr6
yFlRAhbRUVYz6B0aqpLUcf2r5wXDTpnapn3Nyz1FGLYf+vA5kjgFVIQITGOPM5srfTnViCqTNbPL
xmzyXSag+ILncfdWuWHLeQtt7brGKzUdZbCHZPf1hMNqufHq+1ZLu3SmGj3RUkEKg9ZHPcXiMv3g
zZZIFz9ssXEaI7zSnEVdBz720Mx9SB8WgLy6xnIhwRusJiQEmS/fc4zeqz7d7qQxheruuu6eZ9qG
L1st3Tz3yKQaRlFSBwtIBIX8/WJ2lbartJHiv+nvVr1gidF7vxOO3NLQLIzviloLM1MTNpEuWIbm
qUydB2XVOdhuPL7G+XV/6RqeBV4inEb7biS27UaEsLdqZoYkHAYJ/bWZdA0xkkB0gHVNV1vOIrLV
rLHEJItbKDuT/k71YVieAUvKA6d5iHtGzZyixzYYjOK88BZMhEC5bPUIzkfar0kHnLq3MluOurIR
AyNDfA0I/6FxPPfgL7IuYBqw0uOxomBBrjqi8ksFSt9PPRNFeQ+AuYrNHJxzIkCxowo/08I15uQ5
Z20DjAPkPN7iPI7agWYgvB+tUyg73bHALiiXgINik10ERmtI7IFSLvdvLmE6zq5Cq9/XdQ8701hC
KnGNjWqXeA1JlwiCvMwJaJjDOnb6XNf2c7PMlWDnWX5E0Pk8qBD/iwrDoDWSflVhC8qvhLJ7Dvf+
z+qISAKrGnEGPEb0dI8qngZnQ1bWUqB51R4Ii2ROa9KUMHwa0VXFpAqVRUPwvuy76ZD1c49vpqIK
d7OCVa6ngsiX58KBhU//HAXnn31z32Mcdkn19HlPtVlgGRNrddoAiFMNXTZoD4roSbFidqMheiGW
/rkW9e600fhgeRAAsiiSBSk5rPBJVOAfD8IQLGCFNgrNGg2QnXaFbWxMQYnfX60JOikw5o9oJcqg
1+/Wj73RFksrR5GY4KLRJOnxHI0RgJQithqc8xP0O1yQkaJDJ5q93uXrcGGBR8mUmnJHMTvb3SlF
vUpAR5Xy1CbIiWaEqIy61C8386G/x8td9gmmumnCJ3odoKafE4k6hlerA5yK/e0pxrUl4MfqyR6R
ZpAIYQFF5RUFeN/o2BaPVy3664dYZMM7lfIYvsRI1YHsjABNRMR93CQKzVlDYXDMSBCBrW1zjY5z
CmsrmSzyQsHg/beCEfbvUUKxxLlHm2+Q5AtYkyBJ1mvhdC2LXaHsLTirDnXu/IwfT49SyX3ay7DF
F/A6kyzLC74dWaNfnCZztAbArL3aZ1g/PfBSD2XmELe95dKY6MPlCGxgaw27A1jO9n6VG49SIsZL
lmu4nfxbg/k76zuETw9L2IV7VtA7Ayp50nA/PKHqgz7PkqCJq4KXq9gz8wv+kbTG3jSqRuiK0VoM
LTlyEnksMNNtFS82uncOB/rT3GqUK6q152YTTsRMTXirFjZpXH8h5623gqT5BvD2U1LNtQItdwat
+OEoFE3ELoDc7L2XyPSAsvSD+LKVUUbeKqxtKxSSLPcJArLoJgaHKsSHq9PpvyMD5M6bWW9yd9sW
eX5wPVanPtsbV+xNOnO63Dylg8MyFm5HCHktwzrpZt8cPTXEXb+JlCX8qQPurolj9mUHmMsrcvE5
fymfFhcg1CVlCTllX4DLsrGTZ8xC6xR6NAigBqeq/SNtg4T0+vWNAXjYZulIHSosIYbrvyC7U4nk
bmR/BFMLywjgy7vMiCkBEktzjme4OyL0pDYbdn0s8DyMA4x7+ayeNo7zC2+80TuTfheQfe9/IME5
MKlWczV5zjoacm7fII43Szrjmyd8cXLN0p9a+U4u4zSRCMNhXVVIW4hb/TiOyQU44qUvFhRCyVhZ
qLRnG+6tcJMc6GDHcPmoRb2NOakGASDvR6brAh2T5MUAyv9qp1DIXw1YTSYvU2J3KPnrotxptuyH
+KbfGnV/7C2z1u4/7s6Tpm44Xfcs08R8w0kRDHpsJZqsutRFRIo8Y8fglelNoyd82ZrcE4BezaDz
/1gjvc70p3PjevrqVJ2g5FzOp1bLPmS/KKrapUTnLdDwvEDSPmZEyxfnmLkFB0116gCR27w8TO6G
Dl+4CjAC3vIR+gb9oOQgM10jlTJ12xmxsisbgU462FzRqF5afAGOC69/Kv6ngxD/Th52So+EDMmM
ePxi9vtI0UTmROKveFpPIcolmyc69z4oTPmDORLeWW4tC0TrexktNasfRc5CIqnDq+GtNUmkImnD
aElkGvT5INJxVp+z/wBo4GvyPGgQPySb2d0m2LzdQ0I8kzwjo+Au1VfiF28O6s3Lj5pHOq4FRc4u
lOa2Aci0jwKp5eFbo1bKJkYOWfr2/RR1U4hCze6+M8cMyaN+k4xLeKSuR4yk4TXFT+PSWoxU93Ep
Jv3ftUfG6jeBUywGSmtFvxj6UPqfkeI4PGPnfhttmgyokx5WFHuAdOTxEeSbDtOnSAzABPYzsaBw
JG01n3MLlQ73i/AC+VUpSpDPkKjwaZrN2sBj+rujsCH5Dy5x9PVh9jne3CmcZbUYCCD8Jbqhn735
OkSHC/JcqXnQFGMHWzf0Vfzd3NiCIQ6PeUR4hhf2ZN2tDWkAS37BjmfOLUcnTvtW+hMOMZc4OWwI
CCRA3muT5vM7EU87jsU4S/35uMWexXiLBviT355bSX6L85UBGhMcpdN4e24TZugy+OhuR00Am9L5
ORMXhKaLzjEPtB64JRGj4cqMoxUSN4jLv/Kmmp90Z63IJ5dgFgPYrZ8xGSlbTxu2J+PEfZO4ivwN
faxToK1winNfP3ySUM/BbeIRm8hfUlGsGT4Zk/HyNjF31uF51Ztpfx1mEX2CEIF9GhTdRihk8O4w
u2pY1I8pT3WhWjUCTbsaN/7a0qoguY8AAUujoeByj00Wys4S9npWGYzSuPemamrnP8K5rQE2qE7R
FLmYKMzoOVvnvXX90eCVR/7ELCpv19k7bDCCkRnJNgYGAFOawTlhMGFtz1N05lHG+6RQdvqwpAX6
UNFaVYoW+K1EiHW4BOThvo7I2SJmHgVDaLrWwmUo4t31dgaBzHnPC4W4e3Q+brCJMpZYi1KaGk2f
51qQrsQkHUDp3bKndJ+O6k4EOx3NTJNojEQyJAickVAmpCSJYsCz5zbKHQaGJdLIhSTItLKHgiHb
Musj4CANB10lexufne1LIj2gCThh2c5emw+E7qE9I6LY4UAouPzyLNGrAmWy7ZS8YlHg5weHFVug
YZsrHXK+ZSzl1ve6z6fRKreUm/LoPr0LC62Ikl340J+74CULrADv2dO/1EMe2XGbU/uhgzMkM9Vd
0NwX1bP2hkMkTymk4puBDpeatn0mXKdaXpLs+15Mh3whh81g6uKosiwywz/VVq7kM5x4rW99lpTb
behMVz+Bk5YcTIHD2Zp2NwL0cjTxvl9o0C6EDQDBLm8sTBDUlXnjLq3YpIzzsAgIDgUSti4Yvn8t
1MX/hMI9+lplhziDrwQKFnmvdIEg86DHbvP6HwSfptut9S2fp+wqhbMNDOcC1/sTp6OnJZzzyKAd
naI4XJ0YzsaYtTJaUegv2o/+k179OyK4IVueM5aQOYeQx560iuWpYQIkptzgRtnoR1usiTnPztzM
v768wUZhfropzz+LUI5NagtPF0cHbUEUhv1RV1VyEeGt7CrYBWwmsbsSTHXX5YkSlmm/EtJR/dlM
PX/IJCG2F6G2ubu/AsNP6XH1myjrPpdsHwjdSjaWrR7llC4osu3IxKHdm/HovBpPp8xupMwnVrag
rCVPPvdJIOdwmxJQW6dLqMqUb6hx4wSCoI63wUjs7Fb3nqlc9/vOdtHSZlSOkSiWvgUaSPR282rS
IorF7LXra9STv3oihlN+iGVwcZp1HS1PLdwnKXHmCMWwDGbie2GXcSlklQuKUCKEcpgBEoTwIq0Y
bgfH6rY0EA/J4ET6WzLCYXw7NiamjSTlS/vyI0SfotajD3BxqAHq9OTGbj6WANcS53nw4Km+FygZ
zRCIDEUakOBd84JouMnnUtgYQl4SlKQa0mF6O78tASpWV2gFdiHifaVB7GVQ0auIcUf2h4vsIfoV
RrREBM6LUqZDm4ZhY35ZzpjVoRSR3WMXSLsgaUzY0Xrh4/zC78p7/ZNDJzQgtDSPBdXbKRDTuePS
hJuDPUTfW2WjmxbSDJifr8PAHz4f6xLx43wyK3ePMTZJC1LuvUIZFZ6AgODYM2H1Ks0WJ1eFjCiJ
FRA9JwPo8Fh7pvzlFr5wVSZrMufvTR2nJUwoszodVIDyo4RV+eB0hjsXzMymoUL3FUHq4eAj517E
e7Q08v9PeWi7KZEUOk7bddqPKF38q6fTJTf4Qn+hKCsIFvvGyXrs0waq4VnKYsxW3hRyZ5/Z/MXd
zxhn/jtZYUki/hp0fr0caXnrsLG8pFiQoFrw83IjOfzttXH63trxTL6q98oimsPb9diiw1qEwERI
Vqed8AWQ/yc3pNmiCnkuWy/7tr/CBfGLz6gS8TzAtc7nFsd5gvU15Pmb3Bw960yMqxz+pZR2VmwW
0bpUyG6xxgaaPzsvOyVVM+CN79mWuIdsfTDZVoMZR7UNtAEzh7JEil/QS/iaYW/iInTp8n/l77Oe
FrK1IBbAU/wZlzKg6ZXf011j0iA51ITAmsg0oz3EkxJXNEf+XnaxgoAD6g+MLIyTfXqFT64UPfGT
dY3ZSMMN6hzffGeN1h86NjTZvr3lJALIKUCTDSn/tWwQJui0t3BpQITKPW//dX3vZ23br5Yqonts
kmBI1b6fd6uCk683l1HLtOxXG/CQMd4BlSZtHcIqei4p+ZzDSAdpG0nubmUJnKuhxljYwELZbeAQ
hyW2Z62KscfxR+NmuGBt+5azQJB0hdJydcgRMBZqR81mDE5SqWWWTzwO4rvobPMpPwktagRgcdDm
1dEpPHI+UnhmS5+iuV9lVV7X8YJXYxK9UjmwQfOyufC5ysYLgb5NR5IMB0MjvVYcsWNypth+F1Wf
iOuOLF48FhTcxLqAOD1JIQsTHJYHMAgZ/fjBkwk54snh6zJHDcEkf5+Iw1uSG5j2LYFMR0fWEWsq
BE4Cb2r22DgQ0gZNGodcJ7gr5Hmbj8ex/iAfWOC3mFN5XLTyJTSZCoBT3pgkbijN07IsTuZtCZmT
o+Nhk1W9vibzgs7bCdq8JQoFBiLjMajz5Ig+2sCRCihyynbBTyF/poauOXhvyF+CIlswkJj72bFe
7TWSnmhPewk3dZ4Eg8wxQ4FV5rYhGuB+YiMkQusjRxQQgKl1Xe1e0bmM0dxHRRgMl7QaBz+dUrUc
uNkm4OuZI3eYjeQ1DsHc4+s1txh4E4rrwyUTryXH9A2rm4K1QJdQl1f2nIhVb48Fp8J8Y1PDA39b
u1M3NgdBFilQe5Fc6u9qg8NfSylq5/TIJNYxbM4np3DGSPuNk8kVBF8DpJb8LCxzCa9SkJgy/WZ6
4euouTllcKS2vehdIN6sKs7ys6+eOvabeQ0W1ZcVENWaAqPVk2LRbSX7oUIwXzQe4N5h/r/dPM7k
P82B75I7zxjSjBCdhnXrD0GQLmlivfiNOVi/kAA0IvUFleLSK5A5//9gC6dSeyWTEpCg0DbW5rUk
ObQvUoP3hu120JY9/ykiwQRgM7meD4PWNsmEqyWA8NY1+MRMWI3EAERxNHJ2WdKMURlBztv7qe5P
wCSyTs52X478XTZPUSQgFYrJ5lGE7W64WEv6E9uc5u0LjqniqVsABxkT/haas3YgzsTnvvLykpr8
DgphWSfNELYT6TRtrnG+SmJ/39R1n8LdOQ69wOQnYqONfzG5eOfWPBNR+4ac8N5ZHqRrJ1TuMi/g
Q0Ei+prS30QHvo4Jy1l0kRLvbA9rhZcsUN5sXVyM3n7EYAeWYn69aGqN7uLTPsvZTKxpKkne6nKE
U35uMut0zOwfl62YR6hByi4lbNzX3a85FjNQ5w9KJpusr6sWLVDeRrqSzLPh98GGyupXCnuCHYrL
d9WP3OxF8Abbjr4PG8j+1q2TIfFuViXoXKKZfadYqsX1TyFja7LhqA3EuI852MLorKGaoQMrdDhZ
aOH2oC9VMxo0vSoVC9eXxyteoV3cfwG21JkyefZ6fMAzswohTLDnkuCaoXW1YXvLC1S0JSLe1fT+
CKsWTM9WINN0UxGYRVLblneoptSru+6H2dVROqGnZr42vAfA+V0FjsT4ErBdULRsgL90LY/GJUng
cYDNVy40Ie5hiXsOysTB02OVqloeFGn/P5+jriOsE71ZQNqX1MQWbqcx7zSphCuQt+jk72MBXWnC
LuQgcu1WloaaWooY0Ptdjh0oLr0eGg2SBQL3ClyHGBSM8LXxg14q4VBNI2bNvmT7kjctcCXC1r1y
KGvWD0lp7/oTx9Ff/f7Bd3o5bincxEBjV18w32MWhHhTQkKrPOegsj4DQjp/ehJSnQORBBbCnVlS
I3+LWmLfeY29HRlyd7iibdtzlXwKyqjt6+2Cl0Ue8GpAuaQO0O6VF8gZ2HF6rYuVJ9pOVXCwG4/7
Sw9VXuM+0EAes+jFel5GbLbR9HQyqMrg5XpNRUwu5JNAnMtQQvKYilTcC08WXw/tqzaYAnRLnfT8
mBjqzlUZ5OUANYHNe5U/sDkLqzVxu+54BtoSB1vIAvF9xONRCMEfhXGwjnMHJPf0Jk82GqFRFBV7
GPnNRARvx75ng/KbQB/Cn7H6qRkwnvGL5Fifflh/qFBP50zXXYk6PoXJ4Hevi7zhphy6FBQeYjd/
J/1lmHg5Wy1+3wqYW1IYTY4jB+AFIiEf5YtLPjsYEaLTH8Ez13+Xfsgl+X2fIpIabNVBI1XwYoai
MTeMhBGVRB/O77rPM2AdpZGCyVeBEVVgNErbTXAOf+6Xiv0KfhXIxkLn922tmNVZFvGXt2UYvyvq
IZtPq6nbqkINxwL7zuO/rn8uu0qXJvbDsM1FFg9/oHWD5HNrFg+zQPmEKACcbC70329DXOubbPJu
uL3UMCtAWJb1BTAbcZs98NlLPD9MHwPn/TfqmpxRNIhYeXn6CvRgfDJrTzqCrdmCQxBkbU1RhC5p
0CewwD4ZDyfjnjokF4649f9iO6HYceypI9GW+aw/j63ipeTvFYIjBoI0Wy/TsK8qhN2up4KeLz8u
0r8z/g49nKOqadDKnzdk5DWkye4BXnBtee68ex6n3smHQ0ZpcEttswiR3mmk5b/w9zkCJcIZtX4T
jziycjkUixrX01uUjXFRcScukQCNnGwf0clDwD6fQCBcTwVDc7xyj9WU7h83CJwNF+4uRuXBVEUP
Mk4tkJ+u/2oCDyzje8HcWbdljbO5zdC/sRjmJvEl7Im588H+J7JyP770sQ0VdwMHN6GONCZrLoeu
rV7iqTBclSViZ4IYC3xIHMBvOQ14vIBY1R9P3CgU3+uL6aAxTlYeoDb+9WBXZvLbfpqxm9GHYwDA
hCIo0zqoyBztNB23L2flaA2/CQhLFVghk+KNJZ8fGyYxsohBrumXuZsNpO/VwFqEWkDGCT2OmP4D
Ca6VJyh4gD3ms0yCaZuHZINm8jrFCD3TunhZmLdN8B2wCSGeE5uRKVrqw+tMYUYb3IU/ewS6SQsm
laYfaUIzrZmYmn+Ezlzay+JTvYP5Lk512zlzwl0elh04LmkTX+ZXKqyUDDztPajUBMFv1qaY+LfE
3kUAoLMfBUAmy/qPwCVd4pQNuYWRY6/IGNgIY9XCOawVvdZq9BK8hKBeNMVOuot1iuuXBll42NC3
Afw4eSEeSY6xi/zBC9a+GBXtWvmXxW8UA2p/eggFODAYULDjtzQyF5PwNtLINU/3qrvUJ7nN0fWJ
/jJb7VjXrg1ugfhFsJOAClBYQbKkzYa0uGHXKUaIBbZuFsK0YvfYQy11MjAAYFrDIR1R148mQov4
RpJBy1qnNe8/diB+7KV8GazFFYLNjZcO/kWT2FFT9QESjCWqAsNYtqTSx0ygsBdW9qCcD/RfkOtt
QZZOBE+evaV+dR2ut4m4jYM+uH+1mRC8uvxK/xE2s/MrLzrSTE3kFDqOLqHtREFWYxaEpL4j1srq
xlKztGEavIJM3VLfmBDRxDixZrEPucdFdU5SsYtiswHb5d1OSh3DyqV/ndAEZLK1cx2SKSnPMLSY
oYrtXuOfRSBzZsHjtneXPIAo/7Y0EQ1oiQaWW7K0EgaumZzIVl+rtjMzSf78h1JHJV2PhXIRPlvT
c9GbQccXw/0C4/24yN+Ve/XKhjBfplmcTgy527X0K/00B9x4a9Vh4vKIfr70IW6TpJi9ETKNGurD
65M2MXyBYQqDjQhu0Kis8OHkadq0W5ek0lXJpZng8zFxY1OTtnfB5Yv6eCfyckx//H4XJEx/P09K
I6kq91oQYHctGZ7yJFZrynCglVGceg2t8QDrbXl6CvIbZ3OODypjAdxEhbItSdQ7SDwjqpapZ0gS
oJ35ROPDfVKfNgQAFl1OGSRY/YQ2ci64DxlskjSZf179RbtPAKicAmO7tt5S9M+8GG/nbCJlJyGp
SovSgixVzbY+GAE4NFYmhXoDvnTPmWDHnzwvNg2KEKYmESJXSHpWxNq/E+woFkjj05IIq6j5J5p5
m55YbpSqRnoG58VQhzgajYXxUFnJlzO+VimEDrLByMU9JpCYjplh2Oyt/0cOmWROd1kj5/A0h4MQ
eYN0ShGWKaF0+Fgc5VQsuZUvZFN+5tPAEoyFAJPXlkmbMqe98VXYS+7n06UM/kNOFGI1KhUKbbmA
EhrWJeRkvJCIvuRCslbFdNFOZZZb+l8HJO/LN/kguBUNmtGZLlgSOD7dJDc1DiF5EVSEPUvHUYf4
yOJ6Zs+bwMGNNyZnlgzyjTwQzvSmj970rhrYdGIlmcDaJkcMG41GG2B4Fm1iZy2n1Czk9637cEmj
I+F0orW2yie1PSkBP/kjKhNyBW3rOZcykMlqf861UmIcQFbg89eennXKmaoEo6aGduiwzg3fsEep
AtPsswdmblD3lyWxvW9LgpPgXlglFBUo2j92BWQ6RgkbC1TWxpsfdlsmxm/lChTEwqwok2PWoeIW
R2ty1+51Khgf62fATICtRu6Zy0VzY5DFyg/R9+J44kPf6rjG1rW39eORfluI++U3Zk8MnfV8lgAW
s/zhhJNvwTrxrM+XKbB4IeTQR3qu4Kjby31g5BkqEaPI7wo360/KpeIG0g75glTPRL07EcN4/ixh
a1ozK7zYBEODfqJ8hCXVCYSfSGHK5yANPeLm5aj8WRY1hF7n+CmOnzNhVcpnkrFxmpAMlcjk9W7J
7w3qITWplrBhaiadkZnycLOvDAF+3Hzmo+cDYKI/k/mHZwIyC83ht2bOHVEQ3HaiN6QIXqA5Gtju
M51ZEhY693/FKd638++1tq1NOt93vEHiwH3jIrsG5h7IOy9KoQIFqhIn1y8m9tkxABA3XU8FXFz4
akxESYQZLwHLHf6M6/KplFhEcbxridKYYoc+V8LmEJ4t8kvIWQ9FCt3mcRQLUjfOGOHiVK5FqQ8h
cOfZx2BaPC1+GF3oXGpA6Y7SojiLjRLZTv7jerbZ2Er1iZNwfekR+8MJZCc/ykpWbTsb2oGRGFnE
DOujweKDfqfgVZ9+a8/Af+EjToN+H1AbuV1B5evvMKFbnfJRYLlHx1+Ae5JErSRwcwY1mAO244Ud
eza+MHnboncRwdjX3GyTqqmjoKrXp+8F/dE6l3U8PyNovRNxk1rA7cu2dYQ0GGgchQQTfKW3yIWA
s7E6U6ZCKZUUgkjAZUnnM6zBEMeW45o+aKk3jKpp9s9yvfgc5hmA0PIBCw5iKZv9oWrk8bCVxCMr
mEXvarkHSX7Gi7jPbWbUJhvLItOjleuQKqfhGnUYLmZ7i4U7Wj0GEP9kYMMGUmClEU8gWMlRNE1d
JVPUdp8WajGw/ZEa+ekAVxrDXCrYrbIWw9ZFlvKP/2B1YSsq9klQu4YEUOIoANJQizPGQczZNqCJ
jdfLeY5eGEP30QtpzammJxDCu7hXXHXJRYMnUbi8tXlkDDtIqRvAWmAVUwKEFE3KOhvBCe/7+1aT
Zw7LKZs422MJgE7Cuw+zthkGlJSoGtUJdMcwb6zpXKeQGO2t4V3Xo3Wpnzo+CDO5PBdu/sXMypZ6
x4L52OqFCqChWU7HBFeZE9iaDmUmrte6SoQ0IO21JbwaWJBZ3Q4+ZVVEra0c0pcXVfeQU/aDuweR
F2LsiyKOToj+/3Xhg3XWe9jeVQKl9H72FW7cYzDoieBZJn1wUFVigeOMZdGUqtW2Jus3AIxw/IBP
29NRYTrtW235sabNzAXxWRYYTOWr2DQaAsmUn5CkdgO3QdVfCrKv/uVe94VnpE9fTmJhmlOSKsg/
X4Kn8vG/y/u6zrMN7aLAURDOp5g6scqIKGI8eWwIYHQ7547WHo6XoqIpIimrprr5YDB9VhAm04oh
fbcAF8emaEDS4b/Xt83hrerVZSVy1LirHnu9bis3HjRdCstvIQMkECrp+KeADaBlAd7TTbadXqKa
QQbHOH8ZwHJI5MvROJWqROV1ZcuyunYqZcPp+WjNx1JAEwgJYBH+23DFyGKkqHjira3sVnSluI1Y
z81omCfAZTTcOC2UJK1sNj/L+a9l8APiQ7VLAXudsyOVd7rIFZX62lZ1KxMoEvuFEVchFYpNze6f
ZFo6dto91Sb+0gVWx4Km/bt0QFH/fIesA82jLGMB7dtoLqM5CqPBYNc2AW6WLnxCzJSlTKHEERT/
I0axMrZrypyXn2I8g8dENeWORvxe4SzcNLnM0zNbWasJ3rJ5/QApLI15Snk4GPsFNLDrkV6KISPB
f/Z7NNj2swyWs2aib9CaPnB21PEl8uekC0OHWuoPCiCcwj/Wp1dgnkjs4VVdLQQ7pxgsMFQZlR11
czq4J0TdVe6RUWX2ZNy1+uObVMUv/wJOs9kzJDsUQE4AxXAhTrH8a07tv7Vec9Wa76CMu4GSdmr0
V8JLUQoEHE1CjI0u0R+wkvK8cDSmVt6/E5Hz0HYNw81q4vOuNxhjyxsWeAE3lu47+vdb3b1e6oXm
UmKmOCgvzJNedjku/0TRS4PZCWDDFTy02IYvSuzCEdRAqhgkuojECimSf5gQFbmQvy5W78CSf0Xp
+q8dr9cyDKDvZDGcrYuDPQxf5ObnLlwAtIsR1vp1Z+pDM40ldZeSiG6HULA44veXZMbtWPgMeckC
jqFxpuqte79zo67IcC3250DgBBA27B48nvCghi+nIKWYI1L4/4+XktvxNFRljkyUZ6Zu9JQgSVyD
Eg7aNoedomwxWQ3UTMB0JDIxjLd3hAvuzhZ7ZJ2uH/4otxKRqpchgnz8iSglz7gQgUzaxImF62a7
BUwnGy7pH830nAWokVzulqdthhp3ib5TFfovpmroJEQK6EWAtgLiEvhNC4EaLKGn1t7x5P5Bmezd
SsatfGWvY13vVJIUgvFq8R5abeKB2+syu9Fj9YHJwBawlGL7eD7JeROXT1gQlwop4BuNKKyhNZ33
wByR8WipsZfi8ueD24hBVvLZWEP84mpIrlA8Y4GJMlGZ6EyGBxD7ZGlGEpCJmkhvtDqy5FzdiTBr
QZrf2wHPpOuPtMnhMYYHZiyJHiW2Teq5snSm1UQZq8rKyJEyRYC10dU08SpPnpon55/zQOrqv6lK
HNJuB1stSnCAqcowD6wbxTeJ92gaqG+aVNLIvdxJU9/NOx42tKhtPK0T5eC5n0HH0GLrAALy3tlb
EGGPvVoBittJIypZ2WYP0D/9h5c2q0S4VdKTk1XQiPxEIa60DAk5rjdBGbY2itnFALCHSusGIHxn
Q5rtyFR/S3NA/X/g7xipfRj/HJENf95IIJD4rtbiZ0+av25LT+APuayZf0CQ1xG9DfaeRoKpAAhk
rWatQVtD9wqD29tdjT5Vjj+BPMqYdx48/kqe7/owBrf5q+n0gC2E9r52Hvd76Hl9ZbkvFnuHKE7u
jWbrm11IENPIb4Fjg/vEhnB4QehNc+U80PBKBCP6py4ctGTeS/eyI0H0egXb4hZ4xVY6DJcZ2ceJ
VaUz65z/43D0ihWShOqQzuMLyFFOAYvWuV4H0XF1zkTLXSKYPtxvtQtmCwGoJJl5kBVXgZOBvA3V
szdn9eqL7AVHH9be1tovn046SrSC8voVJU0/E6qfBlOX1xVrfmmwbQTjG9fxWcrStsduyWDiylgS
EqDdF4h1Iq8+b/8bTidNWQ34uzgKmYuxz/QM7gJIMB8ApKH8/uRMPyUryhpfexzGqu4wTqNrN6Zo
IGdM6DSB2T0TBqiZZipPMI4LN+YS2/G1fLi61qaCCmx9VQYWRLN8JOQMiNyf0LDQ1SOCxR7H0Dyh
up641fr3nszd+BZLfhTFVeGRfUDnhJNUj3L1AzdCDM1HdIY2OR8OQbfZlxJf6VWwUfoNpkDreUfg
4nHEnzPQpW0TcOwEhiDTRWFbrI52rurlqdyl0iUjmaJgyHrDAtEogk9CarFKrcAT7NXD7Mj6TZ2e
9jaNmLPXaWrj9uO6xNzzxKMLBX3EuTbIryotQAYGzM7eveZx3JVCG+PFqJSxBpRA2BdvnB+SIjXg
f+8gaPNDi6JGgXx2TYLI/qVaVYvSzKAzMNZvL+P8ZBmlV+S37eYFiur8HKSovpgUGE7o/NNFvH6f
fJZvWVropFcKnLpAZts46HnkVZW76/Xl/kja7far5H/sg7/iCL9jndUcNz6AVC5pE/fL7v07pLx+
wGilpNb82S65FzhhAx4o3hGH3riK1KQGEEuDIuEz9sigsBFkFb1xxQcbFp+510sH0KGjOnPWZuFk
S8mByOkK5Q8xH4vRTqQICJlCeoe3XgiuSgdFvAi3yr2MJFRrJNKevn14OIP3ABeThon90DRrA3gG
decGgD0r/bWyFYkxT7UfG9ynIa9dyezujkUA6A4V4n6jk/2uvtJr4Wtldi+pXg0l+BhMqvFs2r/U
IVFUYRbPfl/VGxs1hguN/Tq+cRPIMWlywGIte19eI1X9hjCyj4huX2ZlnPS97Xel8YPPz/lxPCw4
O4247cQuDChuLq6v690dc4HX17p+X2vl5P8AFxVwOlKbd1/NsUZymefEGvdYQFh0LhuJXzKI/oiW
kOIWnnMgY+Da1NSLgaUB3d5nqbx4bK/V8Elg46iTW20MjCe6q1yUEJLx/mILGgjybGfQYsPywlJV
6D311rNbFN2DkJ/u+UCB2unKP0Ymf/OvEwc64HkwWf+LhtkRO74aOoaOYzYGZSaDCijC1Us4wbAn
tekK2fDdczEq/k2aV4Ipb+we5Dhs2Bl6YkguJZn3m3sj/3+mdC+75PYIOrxcUg86P2/Go8POrXgq
DkaepbzIO+GkliyspRfkwr81Trjvg14D9A96Q9bqYy/Y/AowAmAD3sjOYR6K4SCKkSU2QNVp+euV
C2L5EN4O/+cm1XR8ypZ9FTen82omVbHrifNMOHtij2Nk7BjbjE88zEYWYqf+UE5ItS6HrhULmPPY
v7zUI3Tzj8ctZV8HbvWZy/FrC43y+rUU0CMOU5Eyz76M3wl+U6TYj3RNMvfcCsV5tG26clypgMOc
/7afjUwFfLe13iVYZ+++V+HdMHNdSuLBieqytJWk2e+pjYjg74/ZVeevNmYSikKjdUtfKPVzCVtc
GzPPjhUAyjHuf8q1wHBtKIHxISGwYRhcO7cAJboYpu9KQvcBjjKH4t4yNLtt0jtcufFzqpVm0LRK
7AxWC9g3SwvZDPsUt0/qAxvTfNYB/Yzxig8IHo5moAOlTsHu9fQyCEhZei1PmB+Iny/1iCpVrm/g
SWvxiM4mE4mdmpwQpEuU7ZZOKlTMzMefCjLfo5t1sfdaAQqYs1CXaPGSFG0UvHul5FEEKt7ywo0b
pp59xKksimmnYwvW0ikwn8LaTR9caeSWqwGIwKY7UFGuTkfeTBZQ/JmBCkOMjlZiYNpwY9IOazX5
Mg+GtU8qwKaye/PP/Gy3Fy4TjIACtWWHkI7NaNM1BC4k4LvuiNeAYTXYgMaCkrzRuBSp+UJQVek/
jq34CTJtHTBn4FJfx0b7o7ijXPWv0/PdmTokrgrCq9jFSfqSuW0U8VAKXeG4PKZ/vOrLa8ZiF/8A
SDdpqUrMGmbOrSsntZMGTLViDZcKTk2Dzy/Zsys4jh9fSvROGnv4eFz0N8j0AzAE13j5kOiiSceG
Oz47aPpgpHdyFpJBcfMImp7mRHgIsfbTh+lsJM/GvAq9Chy3vEsMCyo8B/v06OEZaQC4fzckV31I
rqMARw9gvrc84Z52itypKTzSc4ubISitHy9FScbZOBGhokuDWFzIrSNFqJrz/dhd8fiaPsh6MwNM
1EeVJaKimT8LB/bS78En8kJ2QLOe/MmkzlKGl9AyGVhWgs8EihtNEbZ99rQMRtY2MqKKib+oDj+v
DBTpczcyUhZ8Wyqe7oAeU97ghc+WXvI0357y9JKztST7YPpeAXoIigOmc/TFMcJhUekcX359C/Ay
VZ/OoO3+fjSg8QLNvhILK60435OzQY2CcJkzGOY0BUQgKJB7U0DWF4WrV14s3vi1+Qyt8Sy2MnHs
gxWsmcR/C02VlZz2VRkIWyGKs5B4QHcORbEddG+VfHmzgQPthwC51Ugu3ClkvF/tWdw7I836PkoT
xHBWAya+frrVHq88T1eds2R+fvK8ZgKJ9xQFbYfgSBKMZiwDNAO6iYqcOHt5T4yKDjhjwJJ2butq
O4lhTmNZxuXxWf6JpnCPbfJZ7JPRcWNPQEXo9Vspb+fCHIqfXwhwzZR4tshYP7zlMOGJMFnioS+b
YViPcZHbmx+I5digMT1ZEAlPa2BOaYso7MlZaQzLG7ME/ocIN2ZnPQX3CrxnJKJ0yD/HzreGDOYu
3amD9EZKFWFciz9S/Qtad8C+4e3Po/iHvS3CgamBfsZnVF6hhYHQamb2X3f4Ce1IFFAmzWh/HKU4
vjzRkhN2Cd9Q7Y5DanygJbhg0ckGYkoCAL5W1dDOS0dUCZ5cDmQA0lDAW6jvQD1S5YPtJcGIQUq0
gSGQZOKGkFlhxvBWBkf7InRRL9kwsGcHEirEjSpsOptCCk8s7U078Sy7d5+Rmh1dTOlyxN3fMMC2
NA5mrFai9e02XDQ3PlsoPeB3BmoYHDRc5wpMw7FYiTsHZfYIQgNX22vqN7XloGBY2YpgPcQwnmwq
NA0ZqWMEQ00HKLhpNpqseSBMj+mTUZ1izd3QzWUU1RLU4eqvSInVZBYT6hLhDhhstDl5to1irhJM
j2QVlPKLfsKnI5jxA61jH5+9/xDHtUq4flAOBebEDGzkAP+K39zZYniaZrM/xsVgUPLDSRJrCnT6
UlxGnw/zoAA4xL2jATkJeWYTP5IbzunVSJXeDAJx2bkUP1+6egP866VCeLntRrGsu2VfWLk/IdRN
AsxRYU/moebdLsi5Gn3b+OSwm5n1vXvBFVCZKCza5aQg79ds9sw6DEtBYSEzISG0/PzI5v/rjemq
XPAZUPp/zYSMPu9XTyq9rzCInypkC/ug83NRmymn//jxhKz0Nu21bF3WDR5AnX9iUP5PHZbT1JBY
WrvouEVbv7QqnJz/4vmFafzVv69WJyQgphrdYSKKo8uTky24Mw3015W+z09cIwyLQ9zE/Y7WV5D1
LFfePyY66EEGWr6cvbe393DZAH78UuqqHz6PmructBBoWDqI5Cr5rwxg9Uq6Y4/I9wH3IUgH4lHV
5je5zCLm6y/z26Y0GEdB0a90Vhcei+kBaVfp3f3z7zDPJ2waTZIU815/oKLEAo72LnQyNBLlngjq
PaYqs0OHdRXByGE2dNqNdAT9U182KV6JC5hfpE8WavozMBKwit6cK46D9DISjbRHduWgsNw0aYKd
l/Dv3RMVBhAMGbA3MofqvmQF9sL07KA3N3Z/nhFOlLfR98wzJSuRxfH4AhsNTizn0pFGsYv7r+QP
bKlq7HJQ1FXNeqaCIaeGotNDq/N4w8jUSYZV7bDnjm6OP4TcSCickVVDFYGV17DfR0fxN/IbfrJ4
xO//3JFjo+jsuD0IMu2wKr8QtiB7EqEVxPyB0F1KCytXsebVrJXgGrd4q+x95YaGYC9yMFh5D4Ix
Z6RWXxhaa655MAQMoPklFw9/nb7eZeFCiB5Oo75lCjiuoYk2kSayYA1NkqMT6kw1b9GMNiaMYUWD
80aOM0NH0R2zmQcujc5fHhsAR9azyUbCI7csLarveNUHDpRggP1MV+do5YWJTpr9flkHEkOGraCb
VGdUYjk3q8zI/+FtOVX3oaYYL9lRCGD4bAObHlTJcaNtXnel+fN4HLJQU2kdouu9gRcVba7/rlKR
lePIQ0zSpo9dd+23PT/rZyXLGjZrfZmWPMhPmx5KQD1V6fmCT/wB+HsLKNN5YkXee3NZKKuVJzf1
+GV0Jdi9JDXv+AS0fTxer8xhr1T3z0mkqj1LXFnz6BZterVKMztDzwrCCqkgtsplN7jAfBx+bALD
KfMRUCKIN/akG9Ia7I5hC//onDE4fqovbqM6Di037C+O1E7XTfd9ZTU5cQoakri2ZwVa49Ggl61v
oOm9rxb3xyOaCuULYoR3Cy6+IkOF8eLmNHB22Co2xZFyR33vUf3chP8VI2R7EF6CmOBPxZ/PAC9j
lAkEHB0wQ0rmrZ7rgF3imtK+LhKeuoC91+RWzv8AJb0Ovw4jJZT+jvKSyWeAMGLz5e0mdla0py5S
UfJqsVUwOiNCr8c53k+jUhN8FpErKZobITOeWI5VaHvo3uqwNqPG7YexUr0AcqnphgWThCd7zdiP
KUYxKPkArArxWqiDYO6n7BXsZ3YRog05N2GKuyUEIDpIWwZDOGzoQ1qhVp98o5PWvPZqyj27EPW8
urPdDzIROVNWwv7lB2qusR4/NtMM9Med9YlTC3V5VY+Egg9OXRf1bSvDT/efv7Q8Jd+ep5CJdptn
PDBbW37XE7+A4ovgoWxZNpSXsD6CJTA8RMnb2zYbgrjRrE69Pi4MC7/EOZgrt/T7rsnrBtyl+q6L
II0jwMoUkEWDT0QpXlounftR0SF+uQzoY5mvCptvWHRWkNoM2n/Ef5/dCaPwblxFQYDVj+vyr4Kx
1uEv5eQxhhthCMxNyZBQnXn8Vu8r4skX5UyXBY/az4NP1+tvDxh9Jg5fo1lmPtEYHUszXfzGDpZk
ml02YSpCOq1QzSr8yrTPbhEUpzcrA6eRuufnGRWglKbN100rwOvUHmgwQnZWlT+rjWlfHB7bE8hN
OEMUDNmIO5YvwkeDhLcLAGC4TFkYh8jXNp4EXi1XuLT7z3CAvt0Dn1BK/olF6pewrM99YmtDsT0V
aXSOdALjfIKF/s/2tlB8L39Mked6hX3Ug4RFosct1R8qNBKx3OsN/dfzlw8ws97fD98V0TCCv4/a
r4rPqTB7K5FjaADZote8QTTticlNLQEnNRV2i1bbRBReGBboouhoJzy6q1CDclOtguIXxMPKoN73
eYNG+BiNEjKidmRPGWIFfnuzPxT0OTcBFUXtTDa0Yl2Oj/Pt14c1634YVSe4tL3caGmJOpWeAnFZ
4rie3LaF5bWNQsxZdi51CO4wC4+0EcRNTIL3ULSUKbFHs8MfdSGxE1Q6sEkumUb5ijeVQqcxjjWK
JMrrZIzTHzJL/Tc2NLL3W9wbJ0Erkk1N0PtE4STQ96MjJiBeI8/6FFBoBPix5nkPJ0XJ8MylVxG7
kOdRE/IUOkcPT5RWV+S/6HQQeHFnK3cIZ7Of0mJZuof1NkVlafWxG5HDClhrLOIQYDKgmnHpj6VB
K8W5PbwRKAWlRSIMktG0bLszzJtHVZpvCzBeH8/c3/Pg15Rum+K1TvxNPnje7IT2UC0ELZolm51E
SQOiOeiB38U7Xyi2Gnc/ZsGnXIXT58eVoPSDhl8oLh+u2DUCGRkHcciXp/PiWP2muSuTBWTKEA+8
EwDBzDHUawz4LPHEmO06IAiOKiHeHWfV+JZVYe8+0jzv5XKZLM/2keDeO4gWNV4l87fVvoBPIQLv
KrT/ncfGrex08H4whZhSQNuTQ2Tp12JuBzADBtMY/EhCUAkDztXeKrOkeFCsTcArRvnbCgjYBmHk
L26yjp6lviU3w8DsYA3+l+a00kWXxYU8BWKjeCHhbnFow2GHDd5KNTeq5AulGscCCinzIc0sWZY/
PpO3PCWQJKEoiUB7pyrOik9EhXIJb6/IiHUJfSUVwb/QlEGnJ0kV8ow11OH/ayfeGIMZs8vUpyAn
5IVcJjK8gYl0AoMdiXxISVpAilZbLerWmK2kueB56qIW9cZR+piC0U318JUp8mc69lKCyS6o6vEP
BZgEC+L0alz3QFjcEmB5kRb7pgXSuvLEEbJqKtABSoj3h6YJsbTZkWwhRnzYa/cgP3kZMQ41+PeR
K2R3T9Js9rumhJQ6GtmvxhO8/aAnfejEvXoxlGOd5I3kpBYUI3ZHZo2JZ4df6hownJJgIe/ITBXf
hAj5y7/VlXMTI8MDoBS9N5CdMNvd2jbpEYuCwKWL7quTGtH9WIp0mgVWUoWaOkZgF0pFORY/4pUF
el78tEd54jAaOwnxiqbYVVvlu2g+VSKTKejjwFyFIR2FoW9DagIMsSXIJW/Z2n+OX5knoCU6XJZR
d3G29CnoKONS84yDcpePU3oROqhZDn8dEAXT4UE/U/4i4l/KhKHXfP06HOXF2UApvr1N6Bdr0FoY
r4nK6cvzzsxjaiAY46ou6U3PxGyvja0jMaxqxIPtDCl1nQQrNJgC6j2por2+tABZF/sg+kDSIXsH
gVgk0fC2XwMvdjz8cWFvVY7Y/5SgUjI1+CHQ1HDJzI6iyfni63f7CtqkV3ocV7vsyO+inpeX3ZdX
Vn450zq0EKTw6KorORbo52XPKPvziCUzkN3yL2pbKX0x0ayNWCYDjq6LQxZn4E7pkqqgcBBKGsbt
7MSTk7lpVPrtDAGOKpQf2gZAIUG3UE0wHCfKpaeWos5yNFDyFM65u2sI2awy13VQorySILy6h25p
u7Hzx91Lz2loBKeKtuX/w8YHfsN/JZtQFYPKAkb8xNun4eHYNwKaq2NoGtrQEtq/2koKkqTgtl+0
Of0CqJ6vVfJNjDMN8WyFEJPfnvGHVBlVLsNEq+BVtyXX4jznhz8/w7jegB/ZCQ3gXDWIHBGsZg2t
qmURoT9Q0psszxD//fbea5bXmEVkb/LFCnNOGp6YeTpuCJP6SVlW9s3QkwtQb6dEHs8vLJB2XuEE
ajnfSpl5Rr9dLeI3U/Jm08zgzF9IKVL5a3rWnKxD433k68wSQQmaWI0pocyR2Nrdn5p7EBy7d4YK
LIOBovjQouRvrVh/h36TS/S4gg3OSP7pCBy9CKOwrJcG4TeP8LT8XkuTaako6p04hfE95PDI+i/w
jyRJZ2MMQZtr3ZBgECgJBW5DVV4gbfuoB7dEkjQIpYI3COehbPK6jeS73p6K/OABW6z0HS3dDZmk
l0Vr2j5RpgD8Vdrbn8oLoFTGaoWyB10Z8wzjAOlJOjuYA52ugoGWxmPGdZaEiWMmeOFw9ARVtCOD
aNCg7eTjUOaK39IXCDV8v3pJFFW+fXJkRjfvaHrMBUnJcJ3tyrRDg/Eh/akVGIQsjl2JBRsXOnNj
HyvR6xOAlQluSLzKaZMUXlJcNntI0pyUaO52+Rgo3BujYZ5rAzKSreBY9JJqaynbjDhsK5tGAjTA
PTb/Y8uTuxc0dF8OtGEjzFguxchj9damOVHNjqnCl70dCD42Vmh68rg5z4DGzxeIoNmc0qMJdmwN
Bj+OM3XyaP4oI5Rovh5X9NojSmfKTuu75XjPtThQMX5dGt5TqphNpkzyQ2U1fqW8Ve8KNwjCUNQI
svcVk2WS6GzRkYtM4N63vMR/e7nYzY+DSlbFmnTrPEe+OrNCjuHtXe/sbC3I/KpNXLhgzMPVzeFx
tjsxNlmeCCNO4hmw1b9QbUD+XeSbrxld+XJFhNaml64MISFHfu+uPctNlEoXsoInqxm7vwSynVaO
D/m/+HWpEKTIUf9q5ZagjWGaF/A92dSWFB04A2irjj7lajMBzyED9/ValgoAZFeg0OP8T3Fs20Wk
eVXXOJI/Tpxuazm3P9q6wHrOIF7H6itrI+bXceB4Urrk+pfWLfAngRm3xFH1rxh6fuaZGsyE5Vl9
83tQTEzd/6GOAXIBYw8CgN5WPJaZHiuIaY9kFgsCY7/BJjGAoHM2giiE8HQnX+J3VUnpDczGy+t7
G8hR4OOQ7fwkM1+ZRw14nNyDPkHZ7I8xgmxJTxMnXcTvuWjK9zFn4xU3tDojlM8b0R0LQ9E07zWY
WR2gDZ1in6xjsmFrBP/5QIU/fvwOABihwRPdCr0SM+MW0J/Ss+FgYWQwqYn6biRmsTQhVIs2n5tK
smzP4wiJ68fWd22ehDtWhgY3ASFlMlhzyERhHr62BCVhaojP/bHBKk1VOnLokxG0YoS8RHF7vL8J
aUWcRe/fboA6yXKcauOvFVh/iSGOUqhfhv9XpKZyOrPzBgDxwivxDkz7JOnpaPPhVRLyU8H0E8wj
h8xHb7vy2UI5Eezif2uQY9c0Zon25XQ8aBZ2VvAd053BT51X7YUitcknZicYRq/IEQlPCcTmTfmG
G2eCxIeFNFCwDsWBlym4TbxiWpD9TePm8hIw0o6GYnAGorde0wqamBLTs8BKc8a8v2Sek96bE9Qx
vJOtZzMv7Pakrlqassj0a1VPpqzvEkA+2nKtG9obBYFToR4XgBodcaUwvrGsPG9E55D2W2WKFw+y
NTZhGk0WJPFTGray89GvBXeEKOMpyUUVD2P3Nnfjflde/I6NXZfIHdwltjDoCiND/DSLiDvJhRbg
dF7nTCLZR4zieGpF2kRU6omf199Nb8CVNB2BLWwQGJ+stTz99EoGPF17uH6rns9BBQQcjhDN+Pak
1WSoEt06qQuBb7lYGPT6QIrbGB9zJjvsUALLJpcpAAHLFnl8LUR6HZo9IoUogDNs8lTFM/Bv+IkT
6uNktWCM5ofSR7spfBJG6gMzzBGtWsdhdGqEFVGoRVgOVkRE+phWD2ZtJ/clU/OjHK6rDLH5pgEd
/BBhyL/i8J/CZQFdpVSESaH2ygA5xJEYouVQ8OFnVECu1rpDndqrn3zQGOeRX6/Yyb2mDCQWxkq2
C34iudmvLxtPW6KrjBBn3H8NaUwkWzwNN+uzvvY0wXNlQnQ08ZZ8M2gjp4lAbrkn7FdX6A4UYvNO
91z2uMePviXkapYdsmeRA4qFLV1ZP5HzoXfNHent2msZposHntdA4s5inoUPNEShpIjLweaPi7Hr
JC1l2ZRVy7KL614ZsP8SkwhlIgpT+ew+eRjxph3cJp8FT9EjJMUkIxgePMw/0G5d5BctWuvHEsD+
8hT3DgzaaVniJAOhvEjjXJxwJoWcLC8pVj2h8m62avUq23PgVLdaSZsyWUD6ToSICME0GpTFnXbu
ZTFqOPcR93qlGnUH3+Upmy/ro5TSKIbKJ19Qvmf8Lpc1qII9SnT+LWwVohbUKQWodjMPgctxpgOw
LErsN1HQfhORVdAmkK+I4yYIy/h0KT6HNywqFUdC/cQaMty6hyGuaOzQy4vICB2gXTEX0jaOUWtG
W0plVSHcvRDbA27X07BGSBnUhtK53zCJHait5YwmqOfdiCHUEQ+cRuMmXiP7RJZT6cY7OPnkx9Lp
75ncJ0O79DUan5B34lqbDH4hgUCMAJGa1slVUoYH6pdyH092PFh4DKFwBrXrQoNZ3YbUDjI9yWlp
vH+te8/cls6cafQalTX4o6p09rgycgULyZ3kKJ2b+sKDQAdffDk2A3/B+1z9i4Xm5uL3mFtVXCBo
Hb5Htb6NvzZaey1NlFnNQVmHGP7xU9ATX4oV8LH/hxauTyGfrUSiceihey0/vaPj0wHxpbAumPS5
TIrzA/SFLvsMC+l8NYLM7/ff+R3nihmrTCWgJ+/fQkSf8C7K+ARGdOBab9TuaTsGJ1L2J+/IEh79
9gYf2JHx5wUgv9OUL3sTSMA8axV6S7gwVRglca9csk8Mz0I904MSTLt0sD3WMexakLsatym4Z19j
tZuIcNWDScF4FCaNj4Z7kbPX07HV1Cj7mb1ZygRmMNLAwZ4ZVIqTbuITrWU8ijP2PLHPhowhZEIu
AsU2oZUoR2poxlO/oUA25NTAe9CKNGioO3FCA3dBJPuCqrhYdS9G5hv23zPYP4aqihg/F3o09Jrz
O/9+Zig2XDqA3pvK2G27mtrcF57EUZ96NxMzlRlD2MC0qL6dXlr7Ynm6ILxZCL+jd1EAMNfeN7Zt
ZIStY1MpGpiE/t9Cr8Bx1v++GS7Q7/M+idrJGrjx1u1F6EuloYXDTUXgqd1sxzUYN0AYV+4xum3c
BEpBKF4UoXUo1mvPU83n2TFG7uWddxUm42Cj8dMFNYZY7nLx87Jk1Mx9oRR0qPAPzNjjK2jlpKdI
qU/gQyRl4oZdVrDMXIy4wtwXXuiXWjsJXZQzV7JhmM6UZj9XZCiwErxZfnFAjk10byWBJOSC1L0A
UehvDG8mzBVYaV9cUiwmDDzkdXFTrfFJoT3S2oltUPJEG1zSoNrasVfKetGxachuOUmVYvfhUELx
QFLLXJ98HE11UuRcYMFL88AvOPkdnuNXoLQiJUwFzfL1FlaN1MGVpoy3ibTfrB1+Z7RYNP1dzcKm
A8L5o1xoTomgyKIW4IU+V2Gi/VaJKTU8fDO1lH3E/CG8cjO1Am3off3R7w3W0YIXFpfVKhHblAG8
vTe+T2293LwQGIHABJdHXX/vNh0bWc0DxynKURoB4DpOGtmZ+1/F7V0HS+Yx6g/p/bqjFXWEp9Tf
ro+LsYntN7SzDnvpY2A+GdL6PVumIn7GhIpqjAEH8OZzI0vn6pWUoODDxvFx4i8TlLVAPjtThP1M
lx9Bo1ikpfjt69a/3+gppuBBthxI+LUqpBnxYXGXIFJqzXewK4SHtRMJu66zhPSA0ljLmmDyC6gc
b6UAblAqS8JN3cI8MWw3VJ0htI562+iOW0451Oc4UjAkmmFo+rQPwg+u/5qCYBnsFMFQNWbw88Kq
FrlbhsOVgMbjDcXOiMMqzBXiKaPb7tU8Ewxb2fUuB2LkmfItwy5euh/SfQw8m4huZ5/0Vsov0Qwl
0BIkU71CJoE0pAek+bf9HybY1gsu3BCnVJMgWta2xvYbv8zEJt+T/br/q/LYd09Na5oUcsm0HGb6
x+wKlJ20ZS0gqytsBF8nHdLrgL5kXZPQvEFZANGYxOgLTrr63E3R/V433hkNRte0xakJmaeiebcm
XJ57OxPYPv2SvnTk9a/LHeqU7hLdTeoNjIZ6sfswYQ4dw/i5o4aOIYvoih+suZ5vU7XwX8WkSUT+
Uahe6y0WGS+ynZc0c6LPnla3yQucw+CIHxLz42iDEKFCQhHRHaiuD7hpukGLUr7YHCFvHsYrAn2S
FlkQVMMOAhlCbijrTZV1AskjMFLsD5Ef9qauj1aBeh2FP2yX75JU2xwKcpgaHnMZbe0rmsrLdg8Y
U2bBdn+ZnA4YphrsxBuHsPYY2Oaw6Q1FG7NPEYGkJE6dkzv+Nj2231aVE/N3iZ7bJM1/PWANA6mD
gAOVSIVm+DKvM4qKQrHMp03VnMMvoCuiIavOgtZBwqY+N7fh7LK9edIgKgJ69SqjystoX7J6uYnz
tQtmhh28nvwP1pYGLFZKhiA0spiOizJsIqhcJF9GXQ+VPSDKeflPsdEwOJQatrFqR5v2zVjyDPbt
gPkWS9k2RAxukzgowTrpbjjG+PcOOHF1MTbhecHTRW85DnbMpBCGJeBa2Tn5jyNQAMkPHsBmBGIH
qbhPOQNDGRXT6XZUP7TbclYKwlMt2+NDrfJPECAK1jPNhoVlTXvYFTM6F/c/xmYS3JB+d8JTsTaH
jWglZWKRDTAZtDkZ30XOOBpYuW/2szdo9JVQ4mnbn1ECJnL9R11bWlVizH37f+FU0KhnjtQfL6sx
WPbX9zgbuBIhceTvGCiAcjGXKsbyK0YrlTw6IgtLNt6l/Z0e3N1zQMxetTwcTTTb/VSqLs2sS2J9
/gWr502b/EP0NHjKzc/DJxmzQhaYSoVwl534bnrByw5UCgaQcqilM68NwRi3L9B5IL30/iB8AUPL
/+TlVfyxSQ1ULCINkuCZ+eRk/02lVzdOFUZQg7/sNzHIR1MRv9Su7YszhsEw8bs+NiZ+nfV5/vmK
WziwPdrLh+dV/xESQilugr8IQwKYUdCiRzHHbj2g9avVJqIR4MfeqLMqR661rgUt1nO150ccH+n8
CCX2EuW3vDnzp9shq//aNPk2TkO5mMMo0qmVw2GO0rWOZINMLulIKTv9E0xHKzDP/fE9XQpNuUc5
SjjlDARbzZ7fWKTaHcR/sbc97Ff/r1FQxgoX6WcTHTsx+olwBVfDvQlUYZFQIBwh9j2h9sIj1U35
IKEsnKpJfNOHwwRAMJeMsuj8lNtWT9ieW1CMCa+TJ5VT4NhJdY/8FPt3TlF+4Vnqk58k1teBV2Hk
ahgLrs0RhAeqlp/SdvhF6HfXLbF5v0RRbOi5PsmL0vNrAq8jxWrObqiM/mYzhjOHStQ1AW+62hDx
OhA8v7kqY8Hx0EcY6n8EjY1Cq5MY+HP2N2nT9AWD5SS0ybk7GXelF8XYAqEtzy3e+cuxAAzU2q/d
Be97sfaJSL6bwvM3W9gGTLblEMKNHqY606TLHVThOgRlVesX+iTynVsl6zqJwZY/hDSY6g2OCOTS
JPmHlxHFOM4o7JfH946QRyTuZLWle1PpBxQUe4RdRhD+xjH3+bif5HWrrj5WTrsvITLuafCa9BiB
QTi647i41Hpsc/MToLPRU6qbCjBu/3wEbq6bchFy0WrcsddWDTRqgZ7tjvVY242UcgR/e3LkWrPp
5MntMWRtxr0WcYkkVgWXA5CnVKcWKk0s88RfjRCTYYaSRCIXqjK8lki4Fk7fYPn8aN1w+YG1/htS
RmVfRbqvajBnolNUOds86PGPn3GTuzo64EnXrA5HMJ4B1ornJhbhyM7DnlFbQT2wcJwEfwbSRE9e
RjuDw+AlqZstrK5uST2bR3yo1n+ptQ46wvV8iDGVEHtPTehVgrkoQ1uMUauJStbJqcBS/N725Ii+
+BvYFNWCsXqUDD+CarvhzLE0+6ArmZC5qNEDK2UZ+aOg7XQLMpGqJojP3OPanXf30fsVeWzFA0ch
cC4ku0iRqyGxoFmGXggQSCTWVoGupMiCt/jkvqF78MOZKT6TRTp86dyZrkWXEHcWsY/ZnEhDHZym
i4FzhdjWQB/FWbN6mjZo7ZWfPCxWN7KBTlizyhT4SMTfbY8DI+Qu7LZLdEU/nmMiHbckbQ3x3ksN
l1s+uyy3TRO3LqVwiv0b6YFsyI2iQhg0z5GTsj47sAydtBTs6AlHq/FHLix5CW9iGKy8cTZAGe9c
qA8P8rvVeoytmaMbT1fNyiIpFZ+thCh8J+ngxvBHiTMpDLjd9KEE9tiJCp5iReylRV5sIoiPRohv
7VHjnqIIz9VNk53xvGooS/Qvir5701s83aion3tndcufQlvjH/HZSk2ZymLSOVAnlcaumTHXS5dB
eIe/koaf7i3ZMZ4jnTI6ofQnDeGhXBEHOAbF2UjJEyfVDvg8vQRN40S0JUJjX/elqa7IGlUj2HBn
4whFS4t/E4NiYEtulJVS1xsSQowNebcEW8VjpwY8pghvwIUCsukA8uinWwmZIJXXh17Nbt/0jYjN
esdmIPQ3sUnCkC0ZFnr6jZI6wTBn9Dsyf9hM1qIBbHyEGLlUdHn2Y/slmLQflFAGlJ079VGi5g9+
R7Dq0LJDMRBFf0eehm7VE4AW5KAe2EP4S3dA1UnmDFRkYCJgv4WozM0uAVjXgLdX944/kHnjqteL
CvxxmFrnPCU1s83v2JZ9VCsSfcv8nwk/UQlbJGCOETH1iYILW26aKgnC0Mauej3r+HCRPZSBfVd0
Keke8dWkdR6xSMmSCwXZR0yi3cg99xGa6LIiuNRr0rHzy8SGhuoNhbLTp+xn2zE/YST1oQhuy6qU
nYlnA3V0ALlOCSWqv0W+9NnbF9PuitrSDfvV4DnRt1i1zpicywXUsr6ZCpbuadEFFjrFU4g1CnAz
6YqXbhJnilh+cq71kgAv+GcbO7XmZ3FiAdbH9otZ8nqXBSBIGUzo3lOTzRbHAlH8rwqD8UN2R8gg
DcCmHuaKBGPDSJ1dkDhQsk1zsOIXICkXyb3y5PsgDgxgdJ2HO5IJ43fYjwH/dXUjjR4E+eRR8nXb
KEtfOwQDU1kcPdl0caCWTzaC/AFhHdqcpzUHEUKdNPxfkyW3jTLMG1ChLTo4QKL8kmm8fHSQj7hU
7xwX+IeQEunotK5u06Gvj463FfELaUMBw53v7O2loAhYZsKftoyoQT7NQD60XH/DqbBZOHpjtUdM
PtVtd1kdIyUu+HAvK6y+9NY9glgeZGIDBbrVx9btzitH2ZE3KxlU6ZOcY6QvZyhNsUEQKYqKtE/d
1WSaYqS18LE5UCxzMfEOhGQBMnA/MajjVadSzGVbI7SQz/o2SQU/QHAER1xL5mWndq+uHmYt9RO8
QgtU1zcFoWGc2bTweFJElE+SfFCLx8FkoTBCKsMYV3/vedVLQf5/fzftUw+Sf2Gd/0N44OvOxVQH
T1Lkw3pYkMjHOsA9v8kUoNUiKLuuMUsfVTMe26O0SoBpgbvdXGARa7F753CzohkUlnB+Yxi0J02i
JRAVz4tljBEibjTA46VIT56mIeDM2xTWHntV++RVDycwIuW1S5bgujmN65pcIcRbyJAL0uoY3HsB
4NtwM5v7gLU2XjcTRhnMU4B8fN3ghbv/8DdirW8k9UPVKU6SPRBGBhDnIxan0m+3Dvn0qB0ghn7C
4swE4B2nb2Igu5+cvRhxaymJzAVrsgNyo+VNVNDg8NVN0ON3OaweK7i55LnZOLVTnP1Fb1aX/43a
36lUheG5PrMNXNVaO2vu3c/xrSjIGT+3IreVMWQhFmFQBPxfVj/0rwsAepGarxic6qChxfQ2tI+d
8GN6w0Aq4s9ODqT/Dzl7KvEzXVwkaA3BA1lTBIt/70gUOA68YvtjIMxf5OaDub1CtKXE0GvMpSh7
eD53G/EB0PNw42YJcBaV/Sh/Ekp3bj9iDEwXa9E4wO4BcDD7aHLG6oQlwQeiFmJxqulQghLNrONd
cpRqJ+E5+m36Bl/JXf2FLrz3i2/nm3UMJG45QJZKyhF+huQrV3g4VPc498cUlMbvaDhQlqJ/ZQjs
oiNan8VhqwBmpj4ocHpV8xi22ZNcwbpydMp3IWhYPaIzgMo5dU2uvgT0N4sPhJfifrTSUxLRZ8hR
dhEHXAmepQjjPSRQH6rMeW4EURlqK8lsR3cZg3NvAbUPKkh6rAz+ku37pvGa5+s7boI3AmSlUd56
QcxJZ2b7oDEb2l8S2xsx5rbZBmnqlAcJCZ4TSfqFCoNY6nz4vgqZR3FhsDCM4KEcjzsQ9w2mmDhY
hIEWfxWRosQ/0ATQhQxDbkSnkKJIgo9oiXwoGy1QIViJHs+PwUNmqJgXZVi6HI4t2eFC2NnOYROo
X2yKDf+K99c/LAB8oMG1HPypMK2DKrz7ywgbOV4SFIZTlklPjbPD4YFZOz2xvpNBNG0kLc1117KN
r4RgG3zbYBDn8wvhFSSJWK+zu8psChUD5pGtVmbjwCUTGmFOAXJHeAlR+dVhZigPsC4+nyQjgKgE
Um2TAlHG+4fFKSGC08denVr37SindDIr4vXzfvLyCxqx5AVUg5yVU0r8XAO4gWi8iuCfcVJqV4Gx
YWNNkp4nSpstcMr4PFf6i27ZuEdGnwcHVHVfQ0qrpEtmUXxredi6bML7OSBrCHmUf8xvbSRSlqC2
LGI/UQOND6ENYmDfFz7fr+RVcJrIHMxy21cLIQixkCLAsDDJON/T6urFzBxyGER7Q0L1D/7ZkJT7
OHSD2QNDqbCUrcMFgBzsIsmDXvw8+jJ565aLwh28ooos3r4wEpL+Pywuc4Gn+jE+t7FTMVAKYPlT
46NK2dSlERWGxdv8A5fJCngSz2CkrfCgwvzSCpKIMtDyfPnR70t+GROBFqX44hR0EBdS3OTq1oUR
0nFXIwnAMAkHqRHLglvUcdWKA/nW1ZqUUn18l86pqBZ2lwdf6nm2tglEI/wubLssXlz/X9nSnQDQ
FAwJW/HdzqYQZIWLiA58CLVo/ttW13JkuUB9y7AGmWzHooM6snm/kf+stdQmCTXatwVWcfWfVJ9W
7jCxI2su7r5fIlmDRLDQQRcgGsol1jKV+qwKFr2U3CadjrvtK4YMAek1oyjYJWkLUr5WEDmxp/p+
quBPbq1BF786wvoVGe4R60ZwERMw3qwBGlPl09wU/NIC7ESwSsqZZLuFyZ1lIMVDA8NrIh662VVG
lLO9xH4fbbXwXzn8vPR6m5WDDBNO8ufAHngw74e3BBSCPpmkK/a9WCBtSE6ZZEr54w/4JmhwlXSa
EMwIoEw1WB7BQkhSrOg/fb7CBuEQUUYzDy5lrrswaNLtYILtwKKj7cc4so9gMancj6sju2YuW6GB
vmLWulDH2/Zth7LrQ4i2PNdkBEisVymy4gxfvsku1BsbKK75C3l+LqPhirdKclofsOGqAHY1IhOB
+GwqYDj6QbiWPMKkRQtL7ixFgetSrJUDZcq/1DSd5NKigkZViALTzrgLfyhHlrWuhp1Sf1nJQmZz
MaCG84OmLxUyZW85QKx5a/TTeElAYEI1dVrU1oMbprpuAvIYpvDCcdIe6jxFb+UqpRhfL4uLWiHG
w2UjfLS+DoU5QDJJIyW6dMIGbK/a5+l/+FSDK0moExkw++i5zR1SPIcC0AlxQrN9fGqIb6U10FLK
LjWOHBKG8yLXcAy70w7LSohEV5e1usfCt8RZHa5gU7JpDE44z4eiYHlB6FuNKc//kPiRVb7WcukQ
skLiHkBLoJlwkYqoRk66NmFuT9ZXxO5KM4loy33H1P9R0dUFneEcjlSjlbHcduANCrQ6VTxDi08I
rvH1urjs7UZaRCsurOFJI1rtRy143CQaWP1ToeBgfIky9QKe3eool5osG5aZnnY9RCcudXEL6Fcw
JflucBTFcq2gtYOh3pdddQE1IWX1BBSwyAO2GUHHDX0yop5F7ty/q9WPacw0kL9r5XH0gOW3MYWS
m5FW8jKf+aUFqsmpQVc50pdLYhbnNemg7n8/4P3AV7gGD1IcvRYf2rjiCIweZk2ByIjq7nivoTI5
XXG+WgpzBviEA4LqofLNe/UVw0V51yHjrTlGVjURoSEypbHSteAXaEOgVBwa/ladHwCQRjlOXXvD
N+6Atd8mV4Gl/hXapGgyV/HnKNZnw7ivqAsBprBF6iZyxD834ZVD7upNCoCOm2/mMP6vmDQIEbtb
Gvn/lSN6+7jZEq3WnuXQ/vF6WW1zWw+uH4qUmM0Uj4MnMYgWepqW3RlIvVeXEmsAPZmkU45BsLJ/
HqvFQW1ZnsLm9LI24K47CG/9lQrDHJlZLz/JzWW718BLg5o2RLAevbG2xDKs8MEDYjA3yFjwi/fd
O6GeMH3IPimpAfmXf59lH0SAq5xY7LAj31Ak3aFbZlfzMB69xrBxlJLuDh9DVPnjBsoa0DN5W4E4
ldhWoDxlzXfKz8tR8+6nFyY1JHzPl4eRFRJyog5JCg3EQ6RVed1AZzhwOCMK1xhwaa2fx8rfeKTr
H5T1ACRwj9gPAjtD5UHE/JqKepg0lhlBQvadQFHWruHqqUdf9XnNbdWOowxDf0YMn8fUUH0XMm0l
+50LG/9J2hTGNvh3ZHuPq/2jHQw9LimN6P1i9N8IU3P3hST/jrWxcTHUTd+wsQQHu1zXOq4sfOud
tQteRCa8bRzB/1ExVv06ldZwSu+O+QHEHeQIJDGhk1Sugmj4a0hvQvh/gMy8u6EsAokjm1ET52o/
ZcsE0NTX3PnHoBDSsrQ3tEvZTu86BpHPJaKXiMoyDPZUhsgR5GO1LWVv7VzIJAhp0YBEE8ZpEXUL
Eud3Gu4OXggB1gcPBy/g35CTRqk2JGTjtzJFiQUKiAzCi2z2fl+guwADrZvmnwfMiAusy2KE7PHS
kkIghN+6w7ARnn5TTpiWSaDlSEn3ZkZUWa3GLA/Dw5IFXDjqRK8us229U4NmEJtd2AEzD/fAAETc
1XHFLpc4Kp6H9NoSvflaQ7VF5e8p3qZo9zKRLmq6RHSGqpSJl9ir/522oE+RledStaM91yY7fsM8
qlJsxXmWupXiGG/wjQ40FjZMQgtZSoLxesT+T9ddUpkZtYKT049X2eLSS2yJe2LW7NAyWtmogHfv
MIuIcKn64e2znnBaUzQUbc9fFj21tUPufRIRuupft7eY09aP6yMAuDwPokVOELb6Vl0hF+WMrdga
gKm/tERMOiA5IA4CuaC/sO1ZK1H0SidsiWrv5kUxK91wjsbMYieID3TDI8k5Tz2IIhuQdVZIyQIZ
hjMpuodaO8oxkXj4DCzBIMIDwGfl0i0M6Yo8lBoWxrWPwzYAZiKwAHXKPtCJ68RdokhW+ELMYwJM
1ieG/RxbQ6qHMlZwkz3SZwuzZnWGx+E8NEreRAwrBHAzferRntwCmRHf6oTCS5/PjLfOEkrJn7Ib
LZCpA0RsC9YU45Oo+2/41fSDgvwZQgRh6sXg/Z+avZcUO7XpyoeSslnwfVfMfuwBRTzHE1nC1ORz
/zIED4rFc0FXlMoAalxVZqDT9bXmgk/JH7VOZmgagEAsJNewSteRqgM4R6iKP7f48Kqc+lwsyCv5
4t0sNVvAXo+OI75VmGmktzydl+zTkvpqPWPeBWHQ4wBN8Jq/RWVg70SboYuDUYBZa/i9uOvpIMtH
WsNhWJpf6KYHWl5z4EkUVDRvEVRW3wn694RWU4gVeBmfHXvvcey3xLGm0mvo6ZgFOpPLZ48ZffOv
imL+AChanLHodcSUP18j78y0Gr+AWwF8s5ZVYqSBTd3SBDwz5yX8I960RcXnH3yJ2ZSCIm6ct2hn
eRkwhU9iZeiDKpmn0nO223qC/YA8Q7gNyxp2Rjk5P2GcshczopWyLKpZ8RB0x8UdQvcwcnJ78dsU
93zDFDS6upNpAbKPTw40MI3tE/g6Dg4d4M8ULNfT4BhrD0HY5YaAM59pTjnEMqqHLq1cgV3h5tUv
Yd61jLu0Cz/9x23UTWKx1JKcO1akqu/dJyjYmdQbdObmo6+AatBV9naHeIilOz3xeOBU44jMF37h
6yaZnJr/nD+I8Uoc9lx4pGZzYP86aAsqE6ZWUu0YxU0tp0aDsupiYVsTFQLuqSBs3Roawu7v3P0O
mP6woVfYnsaIRc7IcOTKyDrB6bCwZtp+SYKZG+EVUj8eAs3MgKPR1J29L7M0ZJmPMhVmCpYYS1Nr
yTVOripJaHiidEtYhz63o3FJwf+bSbgzmr8KZYZtXOQpTM80s1ZrrIzYwnMmctb0z+dQ0FqfySjP
oLp1eVk5lf8buxFyvboCBbKGmwxgrSW4j0emyuGeBjx+krV/e3UUTRZ99LBnrSwITcl6yDCMCa0Q
NGyMcklw54kRYyWC5zJ3pvJdv0eqrUmYf9dx5D9ccQzg6QuQjpDCmLVS8HdGd6FrY242Gq6g5z9O
CCZeTPCTCJzrlt58SLNfzRJTtnw8AtVeOcNJUbfeTqHVKlEV+jMVwCdJnz39UBv6pqNcI/Y4ByQu
2GXLB2xOBs5Dg4t+pdDhXD/SKGoO5y9vxhuklJARMDuvbW6TZfOM6KQyRe2ElEYRL4BVNPZnEgzc
yzAbB5wwpTkZpOSR3LaHK9Df7x2CMvarS5OtCikV0euNqS9xFEtgEG1N4NLCGaOUdeLb4g+9M5w1
XoyU5poTp/D9QxEhXVO4IXvgfifKQUTG7fCYythFoYRJ42Mp7KBd4ao7IArY69apWCn/+/xaMKPC
xkNNZitTONJc8WF4DjPk6lH0xQMYg+kl3Fz95xENv9t9kjC3B+e2vEy34FZyS26G5UGTswZUZ9dI
AalyhoLJraAXYb3Sge/u9CHUMTJWm37frx3gvxDAR2s85UPs8zt74LUiZwxAQRRIAIkj9UyojVGP
nRdT0Qi8MNRNqAxoIWNQrbP6KOX60hQqaF87x+9PdHHG7inb6HMKWIQVTfuX9IczNCckqtW80L2M
LKGK+MMVb9PgI5Yh/jJv+lzeFCyUxIyqrqYd4OYNtu5QYXhrpwgL0xfX1NUAoGyBKReyQzrGul8o
Y3FHlgHhO4Jv8ksfWKNoFLBqdohuarFWDmxD9NNmGpwWF9r/KiF4+Oka9nlhVZWnm2C1LQaGqvws
xJE3402CAFz6rMvevBmV1of22BvySFHThJ8QuLj14OnJ16PF4TCYkxvcqxsHus6NEOUJjQtXIPyc
hdlN16oH8+WpYEK3VT1BWerVy66ayMAn65mqpFLIXgsvQARN6WdsLjTJGpV4OfQNwLkZWdIIpFMh
S5hU6piue4JMeb+4+PChQJMFbzau1hGgFKNQrzlSxd9Rt84eM2bDZvKcNIRNUW6QUSFbEQggm9vp
8J5PTKbOqym1R6w9IjPVPUSRdGtC3fblZa1eoqW5sgg2dQK/wCjXBxkDLuj8wrIhj3FXz8ZVzvWc
xIKkn2I/5DLRrz5CVnMHxRcRecAhTWqCg4RhvCV6koDXu9BLtrxDbPzA2/vcfoWoPpEbXlUKxmVz
Efftfuab5E/gj9D4iJyVRmm/LQk57Si1BblUyABCm6GxG2yIQZbw+Bnp/EQpQ9zD78Lw42JKE13+
+NPr4+FOZI7eH3zfu45eOPwSVhYjxt4scUch2lJ6O/MeMCq/rbXDbIlXT/d3Ak/euiiP6TKgmh1q
Bu/OPecSu4OvSyvgwK5lhntO9ORK4tYrN0oIJ6r+zbVyD8s8yszfCHg1gDe2RyuO87ipChq6eJm8
yyvNMHgMoorpt8SPY97HaePz5ndvqR+rMqBLP0m2V9Bggf70Uj3AHMZf775TOD4DK/ZOQF1jxKlk
8yginb/RBI34LN53nXwFbwuINltnC2Xiy8A0jVNZtDSlNqI6DCVcYm2B+y/Tp6SG0wqRFPAuBRbU
y/+GfCw3S0d8b9EHhf6ZQNYNuIWcExlWpodlOxF3mfSpYv12yS+sbN54fl3LjpaMDSVj48v6lcu/
AceWLEof477VLR+5ME6/Kt0rhVkOnzy/l74dFz+5UaPQg+SEiWL0tUQnKtfeJDObtWNuSNf1qlWe
7ynHFVHl2LcJNm88/VM6B7y+AsHQ6+Dlcqu3SEQkGfi2/rP3sqAjQk7/Vkxptzs6OM6sKawnBMrw
gY0LaDGNma7gzBbf3414lNlkMHgfrYJaFs6VkgMZrbpfYbz2qoqsFwvLLp3RMfC/bjeo8ju1MmI+
HKyJkg3bJb77Xxve/WP6Rc/MeRhKs90iqRZZWdnq03gHQTE15kGt6AE3eTX62V4UMa3Kjs53tJHX
x8VZayaZ6tzfrQQXO0veMvmmkmABndWIz5ypcJxuiA8ymDTk9tvZnzO2nmCE7ZNo3dyxd/7ObqCz
8SjTZzGFmSZuVwkC7mBfmPRxWhhEPvCNXt7NTSPpZcGApdfg2GwExXMCm2icoqStU7pfAXxrmO4U
fashXa6a9CcAb/wc/lgI1HhF8AvsYn683wbzYkfzg4l7posLj40jhGp+wHFRckmJLaFj7Cu9fBy8
PKAova+3Kw+unMsT9RJSosaJlTYXzraCRI0sUlk4ZVB6Qczxj/r10NLkkQDfO8xwjh8G9wAdmlF7
0cl0XXS4nALbbP6nOAzPg/1b6R3xwgzHNRvw/kaXzTogwW8ZOxAjvJ2Pl8ZjF2xL7BG1LOK9nMNb
NI+hcbgC2dT8FsGVkYbzuGS3wdWKIa1NKznMKo+AJq7NrcSrqw4nxsteo7YNHFbZoVWoKdaqAjBn
vZOq1D2c3hDlLb2cLlmG7HFBw0ojNMV7qwIbELIM6CrEZgT4eU6Lx12nEOO6f9Lpc0ff7C1b0Eoi
VCF1ePghmPAge2CabiRYe//GAVDSrvHu4F/r2teW+LdmWS1UWSBC/MKrtXsUbYZ/k4e8fm9XblBT
hoxYRhwzqeJXl6e8pwcV0QuKyNI2KgFI/+ZUYYet/qnAk5U1Io7pdXaigT1G74myHPG3lH3Odka2
/rqEjHMKPPMEa3U5Gp4rsM254xgN4DHiLBR8ln/wvrS31hMA7vqCZITJ+zZW/qaflcVrfZfzrzu0
nZwVi8m1xFb5o8MidNuRKUwGQu/z9Kj2ZuCwayvttoWcs4+K+gWGsRzG06pHtqkI3mnVUkUBDgi7
mHGeyeaCGE5+PmBgPfOMzNUglm71H7A6JWmtO7lnHowhKpmJqojwmXDA0N1drYSacCDx/ivTqMzx
2mOXqUsRN3xoIoayQjr8gZ27LY8T+l4BA0DE3y1KAHQKCWXRlfFxszq9+8LSVXQMcew7c48FXwfn
ExdftNI5ezem/YjEsXZZ4RIcigYLJfuQ290X7mMxJOJFNVJU7yHcKRjllU0fjN6JWCyhugTooR+y
qnOGenr31i5SB4BQRpma3kJ3bAyOTRb7vbX35EbmCDfXYAmPhsapGPZ2193Rb7YSALRVPBUxLiQH
jSLRe/Z7/c8+ETFgjdFG0HYCQwBZw4mrLrPm+NfSD5/8PW6khQn0Td3eweadbtVYleiTxsdOwgTT
idTAHr48Bous8XhVSIBR78DbLQqGveN5NVzNhU4Np1Oet0qgbpxG/nPTNMKAmvtUVJMC8JISd6Ln
s5pFK31QwoHZ3bJYaq7o1SaUGaeDjBxAzCNwzzATg9NtqngZ/IqDQGva1AMamD3q6fUSf5sl0F3t
craps8jgkfhlHzXobEZSi2lcePRAfK2ejV1bgxzAtA0vR/+iXhJashpjj9+g/RXBPRyEcGl0/seF
VHyexNsRFImcWLK5MNDQnsY/a7M8qsewqoks4vhe72hBHYMsswqTH36wLR4SqacYZ0eqSsV1cfDu
TMDlsB0EYkxwS1y+jvR7lbEPv2gPTJAuIVX5Crpv8o+AFCJUhZ6YCLTIGQhbsHv9iBYNHGgU673d
7jyH1cHfXaFRjER3keI7MAit1jvSPadddOTdNNPxuZJpRhqEs8QlQpyhsCJ1JqGbKNg3P1ua9DAS
0fEYMShcFT9PpErK1T/z/PiywLAA5gub34G1zpZk+LrtmIx/Jf9iBZPRI9ZlvKTpTSJHh9DRwB8F
nYrllp4UiXH2MM+Tc5wGFm6QjiG8b1z6kBs1MCi6VzbPhPXLLibEbHZwN0tj3LfA3HmSGJqIFbrJ
Xp6xCw+RiE5C08AT6ptuELsMkYf44NqAZf3PGuk/Mh6gopOLaBUVQkPKdONANxbrE/i5oo0tSyOI
NFWwjrx8DVw2HDYw2OWXl2zLRlT4FtnYUTO1z3IYMHrZqZ8ytjYOqWh5mIbFAoK/TovK8D+FsBAe
mQ441DujiiR1e7Ct0W1PVLitZnouNdJL3GyYIAYTZ+jNtQYbEHnGPD04d5TeA+hc2I86CavGwedg
h863lgnr628wWH5FADyuQUls1zBXufiEJZVZkCv3nwmnxmdIquI+FJCB4U7lGjuu8WSn/4KREfGs
mw7QPHzKJg4ybry+YFZKgWh/JfC59G1ipKvi+SPlCcPDTxYtFJRhL8U9NIyDluVir5aE0w+2XR1w
R/W97TlHYlRdSdJVIjDtdn+2cCw1PAAQ36tJ6GMCT0R418z6qIUTyHXOwfJrnwBFdms82vL/0o6E
7MR+8E5nYNW3eVXvqOjBY8NgjPDeIjhnhvTL4JiOHyBYCHC66tUF6ckNqrTxlN/tOtdeouWichCG
r7/Sm94WMzIliaOdSz09eNCsSDZP3j26QMi/Gz4Y8jTWTt9/j+j/reh/Pl9kU5zQZmgzUZXM7ntt
ha0rDDPMCGpOmsb3cPZ1BuGRbRZrk+yVnq5kAmcRd+X6hvneD3os+mu5ih2d7cp5KV8bBMmHzPd/
u+5j3I39hEW/1dyTNsBrGOkBP8OoN7qP4XV2nADEJVdWw81AIsKlFgu/kJTP/C2fRw7a7ut5YY3r
q7bbptj4JhMjV1K9z+FBID/F2AZynhgZalnKrqGMpXXbt2erhAG2tCmvCBeXYGyBOjxtmh+7KoUV
rtwMm9A3V/eLDwwscB0Jdyu31a4uYfHzXVeF7QQVWbjr24K7EzfwqYpidCfXj4e8MYLD/mkz0lY6
M5NN7221kLv0Ns1fGxQ7aKy+ntOSBf9dZqRHs1ivDRjVNzPWyrOp6GqKmPoXoQwG68VLdIKZlihE
UJDjq3Donr2BGOhr4AQ6zLVEzc5ijTmXHWezkT6ogC2m2Ief+47N8OszMXFP3tj6X3lRY5XTkrGs
TYg/6FS8MyFZ3l8O3hN14eOOLTBzdwKbf9CSdVjLYPN8TBiYlBJYJDG1tA5B/NzZQC65xaTylPBy
sVRfqNgTRYsVFrhV7fzZY24OxSh+zdAsd8eMuYVWM4fGOOFj+ZOIxAbwt/8XhmQWCQ7LUCdB5Nf+
5esiE7O/xVH9n9xzukn3CafMxYRWlk7s9ZszygeU/Nm3L/Ie8tXo2wmrX/LWmP83KAh8XDdIcQs7
C7EGKSMQR3Wyh5lqm/DMX+htr4hd6J5+bnL7QVJfU6laIIdkyg2eSsAIRF/zjM0wpf04di2o8xj+
KvNcMdKwoCKEQdeZFi76k1LhyOkINqbsgdbAFWsakeCwik5WdqP7MGYYhReCvAyq2QADtRoi3Au9
zWgkOe0IcV/5dEVWvuncZNEz0e21BZI+QVe9gtmY9ojH1HyUFCtUo+lt0KaM0x2perTeYqFe9pl0
FGfywaMnhNXkl69njgWrTdoHCFEguYVb1lSaPlbwkiqijBCLE5YMUlxIpkRZR/499hybe8iwG/IW
F/uxip+udZj0NPbEf9aUnXg3RAGHTIBaf//rEXpNIRF39xmM6Pj99ySejSt1Hc4ZFVSswS3NccqE
Fwr5567l4klhGGrH/N5pH450Z/dP1DhKLKlua2bMo2DZPV5jpGtIVOqId/hse1onEkE20cKWmIo7
HDZ1SvAHjtXcu+IN6jxtSHZ7EzwA1K7CsbpONqPxoBqMGRgzMv1F8f66z1wrphOGjTPYxqukzZ2I
poKZRO7E7AwesIlWFGUrFLT+VCpXm03mT7rlZvW2RZ67s5VsgGOH93x98OLsUzOO3viuAsP/Wv6f
nHWG2iHc56JYTyQ/tGZsYyH0hsI8dJdx9KZk+aSbfmPTD89CuJMMpeA98I+pslf6ncmlcTvki0y6
n9GHWk0UB/608+Kt0b3ph9XFDTqCLaaKSEaGs5QuI0O3Dw5nfhDs+k8V5QMNsYFVMeajdeIoa3a0
oXn/bNO8XVt2kRMXNlvsqhuPAqxBZqr5g9h0DH5S3q3uEyep9BpB/lCPqSa8Aqc+dzTc/N3H1qat
HYKal2CXX+FTTBdvpfkLDOwdvEvGF07C/lWXGKKupJDkd5TlrplYQnH83U3ni3JfHQssyaAnIB7j
PcEpHgfEcKtT110oXNfvtxABUZ3SiYrUVj1xWDKelzRDvSWyxLfabMLuRDbeJm6XD7i+xZv5OsqR
vEe3GIRfAgErsarUavWQIF0QOKJdObo3v5ztHREU8t8FMsK03MbAqTG6o3lpXuuEXX9KDRrNO//e
L0hV/bBVx8mXo1h2ftCmHhHzHkJXPo+ldidoEOgpPgEa8OZGutOpu55evGDxkHM005h1WydFrmoz
70mLPyKg0ZJMGmgikzTw5s+Ov+idM2dmYiq29C5khNturg0hUyae2duuU0mge25VVWbLVOvSIGLh
VlCr6TrkGuM4dOHSnW22YYfQZlLmWBvZeSn2XJmFF0QYYhBRWEfPZmrt8Rm3OHSmk3qnn2slcL7F
VCSYAIIWLnTYlVSI991ewr5WbkaTWiqeYWApBIx+nlG7V2KKmuNS0DZ7tGgrdMPA0tgAdj3FaFjM
lyzAxUvjUnk1eu+tYO67RdrTtEkLcplfN8HiNlrYNCPvqxrNfyO4eC6YDMYLOTca/JuB3hNAP3RD
K7a7vl2tNXNtB5Rn5LfiTVSqCyzzjolOPRSOo6Y7OhlN7OWkv0/L68J0DTvZ+fVd1BP4MYO6Jr2T
cdLhkf9gfqIrYVGlMxx1x0NOoe6LWpw5+8/i2zeZ+6KUdhnbqqa9DRMsmOFHBevHtWNGTkptt9Er
kaMQNU9hOSu7nXdPYU3BZQiNXx8xJl8MCCozLGwYNdLsJeJXzNHQe81Xfghs94jqBA4PiaVesmJ3
bNfyMxa8RCgwHMs7yOMDix8/iTHR5YCOfUfR3lOYtP39YKY8hAkTlH1Os00NAAXMLMD6VVg/7Yp1
LW8ko2PB3ONMlv8hGJ6uL5KMChrKZDYXqmr+I0yRCrYmK9n3Z9WuYBOpIXlM5ULOAY1WlOoB9UbJ
FzzVW6JCKSBztDLP8Si0rIU7UMGbVvLPFOh2YOyu6w4XA5e3Z92M4bKw/wgPzbVbPr2mJQ6IOzoD
b0tagmN9vmgUdOtZdM5dTsdBcvulx+BXd4cuGp3u7wITv3QoerIOWcxkceY7eJN0vPMnVrHwJf1y
g/SzceM80hktquguPArV5OZ0ySKGrw/5c1K3dW8R1wvxqrylvNedtAURy2Xfl/wCxuCCo7JUQfjQ
w+lNa0nGyNybnUsUtC8GOhIDVFyqoPokdPgjgfg2PeTotG79PcE+c2Bf+MNtdIEtCeZAgbCAHe1f
X+V8rcVIWkyM6gRFOVCGPMMfMVa833V4IzjP7FUDVvyL/peqVvwUi55VNrva8amAm/7ECoNHjTJc
YU+SQiQEcSV4zLevz4uhuJHX8AGrIe5IUpwuu71FqGkWDy+EiUzUhRe/Q6SSEK5RhjvuAyhPaAom
+SrdzHi/9PJCAQk6xcIYKp5G4S7TF2VrsJzn/Cf0GoWZXLrFEbhy0O4az0zZE2EHqHKExocbkbec
WmmZcnA51FdSYhTeJPULAUmU5ujxQAW9/hOGrfCipo8Po8ecvy6c+MPQFeZ9noCiuMyAjselu+Ah
t/H2ImWkdON65VXnlJP4keqYMweAyTnUIt8nS0AzWPOBECjcF9VaqNcDoRHmw99/uW2wZ75yGkXr
qsj+Q8cHe6cfU3+NIS+Qi7t+TDjpd1K35nwL+CMHpivyjdv7hMzpiqSsmdJkCdbpb65bSZB4Tqo5
waTuxsmA6Bi20dzAJG5GRTRrrLDLfML7Cbg8km0O+dKpLuqQSuH+USFt5G10dRcAuIWzap11tiQ9
5P5Q1B3oPn+oArDZhQkZC5wpzreMLa9sD6AY+p9zV1k6rUrjqQkG5EUmVtGsHujMykudDmWNVQlA
bGJ6dZo80HnT9LCP9mx4k4UG6h7jgrO9kziv4GLFN4bwyEuwet7uXzs9YQex9Ra4l9QxQ6B1Bq4L
wHoEh02Yr0EAd7/HmQ8P3rIkgcuJnn74VN4QCgOfJqY2QJ/YCQm/IIHuUNBynmE1G/MlFy8vQ4J/
Vb2etmN8WbrpvyMoHOWlIBBIboG/3r8/fXriARJaYVhh0LKwwsUx4r4X86NtfNiM27iefFkdEFWW
R9gVfreOoeF9poNiLITuz9C8LpMStcTAUjVfIYl5Lo/H0T1U+cbR0TXaIRc6t6RyoozY9ER7+DcM
PexvIx9y5O6RQYHzR5RcTymXX37LFBehPg/EciooP2fYrwwyCpFYb7DHtaLQwjOXFbETdjvH9hJE
e2R2HK9FASI5A+wShCuKeYrw13NwxpzoWGNHqkeQYHF4j+jY1XPOuSK+DLLCIH00Vm6I0e4lmx+s
hDNjxe/3cli6S/9wFfPD6EfzXxSJFhSG7cshDj+VzFs8tjMAblKGiawZNjh9EZdXc2BqeHSZxqKO
FIZgOttK55z/r7rq8ghKiKcwEVmpiQzMRFhuzYUokpJ5DNZmxbfnZQn1fJ379r0LGREWCPrv3Jaa
oRKbzPeVTVZ2Hp0xBGUe/ZubU/1GyzC6ei4FSED0QOmOIywG7qtaQNCf8kDOh+5dbSFYVzBdt/Ze
abH70Gktym9v2Q3AlI3A0YSyJ3V6JoTHEJ/Q6fXpRyI3PQTvlzLTXbIhhr5/3Q0N3LM6r5IvUAgl
1SVX8QxNLpL/hTIJjkmvq+P0wDPkS6wQkmSzycHXVf6FAbOuhUQu0XIr696qshJKivGDosPVrebM
9wNZYqg4aTkFlQcQAcveGecb86kB5qtRVHGyxy7R7/BWuiTNH2H+/vX5cYAUa0ugaZs919u1fsvY
98A1FnL1nr6AwtKF0sIqqqzQ+40jleiW4FaVNDvZpZ37EPwx8IhWQ0/cBfFZffI0OElv/NiePdal
txYH9nttPel2jVYXdI6MbpvYb0ZmjZCEkUzpBWRL98hWE7jSrvm5XOyhymNzXBnjPD0PZLJb24Ya
tDp4YNQ/+/KHGJOJ7fsa0dCCVYDFzURur/ToZPjmdYi7YCcrCAIKu7d2PrV6UWDlLK4x+/ej2agj
oFiuvuwJz4zMxr2zfTv/a+edajnAtSgaF69NCJV7vJQY9c9eOCjsFcFY5fBmjmTzfOFKAvrYEy3V
mQd2IKu9Fkd+1/0hdn4NtmgQCSzqq5uPciu24YAsZiMLp33kKTu1FeI3ChfFjhsc5gnRkdKBWw3c
9pGpDGxFQKKu3OGXsZsrzDeLruE+vUHveKP1WpDvhePiXY0lqe7kUbpIeoH7JpRvuGpY0qNjDtF+
fcKF6uZHxbSGvxmTLWFo7imq02fRYF40PQTQxFT1ucE5JSXrQc8UnMtm1u/07Cj4G7Iny4q+CKpF
MIeXXhUjp7U0Hz4f+F2gN7UaOOMzvWi6kIxU4CprBdJjxG9oMHgWz2RfXe+77bb/tMxnE9lCNh0B
0ElVHLg1fSG/bOpBXdR6+qNWFt0DmnvrG1gM04AmcPEg7Lx0kLfhml/hYB3AOzEcK81p44mrAKpP
5P4Qv2kdu/osxKIWOr6BCnnqRntKnlR0P2AwnHmk++elI2ZJa8KAL3PfGzq3d7DijeBOEbQfAXvt
M7Y+lyKJSNd4iFZ7c6QzFa0I2axiYzRAnB1+NDDRIf63XInt4zO9PZqqvEq9LdTvamdAcx8XbwAJ
5PeR97sZ2bJ3JJCHiBkd9eqWkeb7PaFB5McupzNGBHnIx6dyvGUMO/gtXMxJ3NAPjwgPr50znTQx
Ld5BG8Bv5ykG/lC1df/uX52/qA+++GvDpxNMw2Brut3nKdd77yV8JVN1JyTJh731ZLnGPdicfXPP
st3JMXyIXq6TlK20nqyo9jyZibPRtHEwKhulsFPsnqnHOHNc0JJ/MUnC81LAS60NWLLk2D+U77vV
/RvBP9uLb2JMqQvItD1z/m43D9wWIC5TG3vr5LziH9IXGQYBbdv3ewlojAPgwWikJGhv8meMXn+Y
ucVyqGnDL0EK0Fd6PoxV6ZH8zZKC5wSg1S4bKzibxsn1XtrtDeU++QXciymP+MeNq9zKOtIerS9X
Xol+sZMHuvRpF60qpuBEGRswEZA+ylBkenld8ilKzggk+P8f/i3VQlHqASR/OunuaKfQ/un37y57
iAc8rb5zsGXfOCvLwOP/loHZNfFdPWbXa4cpYTDbHUV3v3wBmBNZ5QmBn6HtToW4297q7LATo38v
rrwoV5e/imW2GVPw/OM1283ddbxyTfCDRh+iz9e1iMJi9xASdJ0MJYFaJc9Dg4aWBn1u1oD6EATK
hOk1FoAQE3LNP3ag8EKoSLCc3clIkN9QDb797vcBrjPE5P3Y0rS9s2uegMeOOWVmFQAvrKxyNyyA
JrseZwOqu+EghT9639OESl2ATHQGNR32Ip4P40ILYD5vCuhQLEhcj5rhY6aNKKLAlPU5h3fWxzAG
2uuLPv0gL2MvHh5dkIRPI3MIh9oD6UW1avtX+fnU4X+trauwCltnznAI1L1xbg5UNZSG9KtYadME
5Q3+B36uobYlnQjYxxI/6YHCQBsBR3xMnGtvgbxG2UNZhvLPDOubn/0Zrz/c0E9xB4Qm0Ubd7RoK
Zw9cmL9nAFp8DPSqzGZf/8o7NIwNSWn73gv3z+1gSZJ1Ch0sPlTHvpxSELFX27vQiXXYPIYqSlld
996AJOHypURm0HjHXd9MM6foyldGRIbkVEfgADB0WBTy7yMpC6lgwsT7kChQZifyQT+ePlXvHrTV
fFcQi/LJzGYaN0dySBDr+t8Du7LjdZvfeWqGccEmA7V0C+99OImFDYiSzu5nHMMvjE0Yv178UFs0
NfMGX60EXGoLDzbhu0mguvxnvFUOEFmr8ipK+/HzVKT7RNGSCl98d1ZPOGrXk7C+1MIwb+wfO6LJ
cNAfKtdAlUzqyrxQaHOcrzwAe1jLEvWKePEMICxHZXTPfpGDJ3xPsL89DMZKBWXbBrCu5RiDnODP
HovdPLjvf7c2if03k2I90wm+dMlgUjcZym8L/e//2ih++6bMZM7BOHXT/kPINgJeYUJF1Xin3Z34
4RUVIp0fQmNRLEBeZ+D77m66XlF14q8bEwoCeyVVtSVedZhr9jjJrlTuMOTGc1KInXX78uhw/gJm
/9K4VEhSYJGTLSYdAZPRw2jhm16zSNk5KVphZq123i8bSZzhYcSdvUbuC5fnoiiNeO5nzNFMwWAK
gPZSTN7hVYFHC1+mL21TcCwxNwmQfMX40ScCoeTC3D4s+5N/0xbtWckaStWQXTbndkvI6YidtboS
3WY3K+PO/qJ2TFjlUgodhJR59/MJF2t3AJHN3GyFQw76Gu3e31fTM4zn8OO4HptGIGIlgfM1WKtf
oMm/SJpSywhenH5K+EW4wm7+Q0CwUB3AOHdXqLuQ0Ci5DLLLp0ownXE2DeyYY9ej84FDbYtn0j4o
dpvsHhtuZFWJNndf9PPpsB7AQMPBNKw5X204yFO1Gz90mBR2fXoli9lOocAZIq2vLA0BX1XLT5m5
aXk8J3vko6ZGsUOFuxDgkS/BQb1txmgp0aeVNpkCz2At5d4EhBtHszdbcgslP5Ik6JDTcBzvDUpD
g4zZ2gTIzYe6Nhu4MsjrXofMIBK99TBIM4UL8t5SxZN40+ZgctaJef44wyPbgMZw3d1QQe4nnTtz
VLJksnPSU12FzI/ATRs+uQDtWLNDgP9XTbdeWXjZAkbQPY06tIpHbcQmLTdvWTFbhbOr8vo/kv69
AoCNHkQZmbSJUteykl+bwKu/EkyNZ2lY2ODXTQ2x49g2UL7qJtAx4a1UF4Il0agBQ5gxRJSJpulr
CkfmvlkqJNU4TD9iFQE8mEb2AvE4KzkaXqUJocNpTNJcWfMM6zGmGMOktOKIDSr3E5zYTNusoaZ+
GzdBziySebdo7YXt5RFEw33jwweRmJPPykiG8VSPBtIU0+HFZ+LcrMqeNke/45UYUyYupAKEnEuT
uDGVOrLeF4YOn2vqMgzinoQaxxyis7QsJkVpRnXpAG+iz+bjOQAlwEXuDlEZH4XZ7WA0TNJ/WaFH
sWa166gMDV2SsfXsmwh+5hDIRS8jcC8rDjO7pTspADYkTmfLw9MIEBiExrQ+KVAk79tlTGUW09BX
xUsPPkmrITbD/x0v0jl/kQIw9tcSM8WjlJWAXIMWMZfrbqfPq9q1OyW7x91/dzaRYHXzh5mlNXRG
1aoV13lHUHcO7gqVOICeguen4TxeCq1rkuCzFmKfZ3dnfCEI1uvRlpf3CkTeolRh/WbB4JTXrzcy
P3WNIaNZFiqWP2kGhcV0NM7uH5d9Y/JO0phjBRXT9hUAsFaf/s0PhIJyMXHOLM+uu5KN7zU8iUNs
JX4HqGW25PI9v+gq+CvwMsulbFhW126trLTUUmofJ/mwIy07CQoqQ4jrA4UTXubhhN16dTkUxudU
0DEuOKDz9frnMs3m7BRzkyZU7QG+m8NoQHb84Ue5Yi6XctQp4Esx6TbAPyskhTSM0wvXccyn4/Kv
iCSHtisbdlLdkYwC1QWcxymh8+t9BsRrVp0EWZAOS9JfgzkBYp0E9g4Ysf0X9ZbN/LK+wWc6ym1T
5qQ/bVvJGNTduFoRRx36qU2S5dWdD1bZgNId7F4yQmxN+bRtm//fv+6R8RpCMlM3ReAgGwU1PvYq
q4vhxvC/zvz+RZU/19sic8zMP2bBdTof44WaEKkdlMI9choWZrjaltlCH0VuNBgC1LfuAvxzvhV2
Bpzgl6M+F8FXR7NHnyZKKYEqdXEJnqERDqCh6bZtuOXIBBEhKehms0KamqJqTgV70l70V3b8De69
RKo7/mmQxDE1P6M311vXKOUdC37GAs9SgWRCYBc4XKGYc9GXMbpHgo8k4wlWtIYHNLaL7hpb0+2g
lAXZWYD6xc1hvbPCYumBxyvad+NKpljxWmxV3RyjAc/57/1ZIhJ5beU0M0piFm7pZU+Jnrmv3JIg
a2jIb+cPsqSoQq0Bzbze3WaWrQO6Yte7NLDu0+8A+85HhWsdQjJQkL7gaKcTM5yNWUADqK5qxwx7
fJhw9qIsGaHK/O4jgfYVFkIr1Q2Xdxz5kW+ovWFOuUrLIzbe2OCpTHkmZQN/7xhAyMsSytFTeNLC
m/OVYrxRJz9k6HbX78H8sDtHA8uWqQsVYeaPwrC1P3DmKU1yYhmtN+9S4vdgBqQannsTQLqAwcPQ
71zRp62bLiAEP3/ACty7xBxqncQwSJSF3B6sTMJfmTvnuqJbk2ddFaOzOW3qFZXJKx+zA/hzHpDJ
OrkHLAa5MTqd+9i6LPVE5V5PWU8pl+r0W+qtTH2imMUF2Q2JELY8tReufUogiK0voRckRv+L7hQB
hl+7bBbdHgNsAaPDR9BQZbbB7ckjLF5Lfa7PLWrsfQ2Kta0Rmx47LwGnPq6aku8jxuo4Cct6F1VW
oXK9J7nnC3Y6leyIfQIblf6zzOHGuvDbk+GnNWj/jPJIEJ1H8UfpucG/YT6GuMGffFGbZHcILcx2
Stv1xaUIfrrOU+jeu2VF21YyXETaIx4UmUWVZZmPM69Y4YvphuD/lHLuOqReyzVnzsFiq8BQnBGI
Xop7fqB5wf4+Ix7J966X1DzDP6Jz+zM4YXwZx8OjaxzO84IbReobQLz9D92L97iSwBB+wNy+jQVV
EbXQW3mOC56uk/b2rh6HuCISfPVBdguPwOUvXXXvv9NFH3wE8c2ihJRpWw3d5ht/V7LmTQK/8U1S
bDKz47Z5V8YCbRoEDhMwzN6n+lGzEeEQPBh1tKIhd/4P8qbcUV4wwxuGMd4e5yGLwdygYbEWDplw
fbWXE/mhN36rwu2JobUFod0WrxI4Zox2pGqBuz0VB0faVXvjqgq07BlyqksLIy3qUbLWn7KMqqKP
Rx5pufPVpWP3qLAatybk2it+oB7cgfAZ7rXNPiggXEH5IjEGIMaZk5LQONCK4+GWFGMUikEcc7NV
TZ1y0g2RUI36NSNyYF8ly/fmOo9yhavbgW4dFLfa+BX/BlHWN+969pHEKLx4xV3GRy+402vbs2ce
xCA7ZSvnts9OqNNAQGOy0EcDAv7XjTjmGDeQi1DgsSjVEBHYVB/tntLuVxYhLhPSKV5wNQ3tQfMA
pC796XUSXNMFwBUnO6TCaeQohpoVH8ikmPT8hfYy1P5vPrzvkisJUK5JuFs5onQboj/TYmOe+FP+
d9UTBpdhGd2Sk0Xyr1JcO6Lta5PLshF9wNWm/l+7IfhUh85haaz46F8KN52pUg18gqvoSMFYfIvN
rHs9b1LjUDNm6q860tjACfN5OGQ0MM54m/7ykaJAn4Ket1kcPpzaXzrm/+kjF1N3SAFcLnHHmnqZ
vLuZLaRfuYqfN6LXrVW7yejQcluATx+H5IHBJG5uDxJAAvDTxzW5TEE26gO1Q5EoK9oClISKkO29
BSJF/2x6JyBoCd+sppHcAVGg8v0xTWBeu9elIW84u2+VwaYZBwHTaUe0KPRT5CPwRTV5dXWICjZg
XiJeX+9HdbCWoOrS71U7lnQJuzXWzNVEnEa1sZIY7eLtAwBuyjdexqyGJfUV2rEHD9cdV6hYSx9E
HU8oGDJgebnbW715d13gGziHUKqxO86mgcnsySYIc2QDi3tHsVxSd+EKNIHLH2T5FKDXDfW6l6w7
yGWS+tnaMWy0fXfgcW+DVkc7BrTMnKtqeUFLO/6cR4ewvOtAkZIsHNmrsJu1Glgw0DDWvkAn/T1Y
Ze2en4p4N8u999QGS/D3bwUY7GlB5vbtMyc7LVK04yjyOGPEudP8izJCeQuCBxOsAqoMQ1hMqPMx
HX4hynNVQk7ao1oiPUVht7+hnJXtN0ix0GyhT7C+uOCCBu0swmtzARTGKfqJR3aMwtLnHFWm5Wyr
OMRjnuxpKbivfJ9FckPde/vcII1apCyyfEKWjHHKYCxNODgajXmyjsZklMcihh9vHi5W5epGh6uK
WMGyB4fyrqahIGRFTrvENg6P+4eKbx1lXoekTGQ+L/brRM9CkDw6fn3JAyJBZGIDxLfJSJS7rrZT
ZYQ21uhZfKXJJDLhe7pmc03CG60tZLY2DycrmdArdOt9W5Sha9opIUXYw2VYnHPhRojIZE8Gc6C/
a/ThWn11YGPARdyM3wiTscbkPhu0mXm+taPSOgUvYJL+sXTMgzUIMP2xv49VjUvS4XbqQ73zZdqI
yGxXKe+HNS6weNw1WJ9lOR149vtxQP/KZjnkEhldqANvbsRCRn+VOypvnuvknJ/l3kTgJdJgWbXL
g3F2MISuHmhRJupFIy30IZ+5ZBkOMqMObGn6yrv3Ljx/NzkWblAYrjqwiJ1s0+/St6Pndcew7PqV
/pDm5aQr8ubuE2oea9rukU6ZZ0ad+rZ0tUyCTR1XF7WydZYqaoIAtF3u0hAB+ZjbltlvSC98Qgk6
NRmNzt9WkYRP9BxZJJJOS1Tynw6q2cBsBxoWy/rRFTRcpUCyar0VUAD7Ih/gM/Fl2Uy4x3Cnslpg
bdV27MfKC5puVhiCSvG1+aetjXK9s6Rbp9cblKJrJLU/6r5Eh0e0h/uXjNNL8TaRKVwYuO7ph60q
ngiRboaIbd3Xkgea7qMgLHGi0q4jPaQt2r5Gr3pM/D3TYw1LGfpH9I5/rn243L4yElsV3Er35sZo
qvIdOv3EaRWWxpe0rXfa16z/BoPO54fzyBSllWbOd7BVEtyVNYdo19T76SAtz9VWmiZ3OLb74gZ0
gqOa2PSnazAFMIxMmETETT2ypiSOapIU/6NFM+0hslhaPtHFWQlbPD1tHv5Mm2JRgsTh4km4AWbp
MQ5F4WJrfN81bfoyMBvITvH4SZZ8MuUXdlnmTxED+omW1HuLca7MX+3CEkA9/RQ6MPqavA5U13Yx
CqzcRGW4pAeNALHLwTO3JT9B6TtfcA/ac8KYcUppAUjMHeCWVzr9nv9NYjANzswtigL/ziV++28X
tPfHb1LMMhhvwvsyecGybljGsSoksvGhbCf+mXy8ZnedrPugbf1CVh2Ml0JuuKNFi1zbp8r36da9
saBqzDAaFZd3EdCts4fIkdXDAFlFjahHLISy4n73Rh9LW+KaXfBUItT2HIXZCR/5h3WkL1phSzVs
YBXQfZszyFfssKZOeXhQNwjBaUOmQfb98osxsFFkF2RGdUaoswuxgTegUhsjtVdChuQqhDM8GNRz
JTNbYvbFa+DQ+QbQ8C+JUBHgfNFDpKe4KtqeQUeAxOA+9mTdERCCLD6MazMgHbZ5CVrHrhPEGBPH
WuGoQ/b5mNwFOcwrgI8a0yXK67+LOf0xMmrpPN99TVtYcl73G3AFf+GpQR174x2EVJvUJ5I+hQRc
6lkn9hrc65FxzsSrbRtP3/ke7ibk2GBGyWoS2trsNYLJ27l6lUZHJoqygegh/0RtkH0H8j/iD/fk
c1PIvkF4jYC/K16NBT/SYXznLrUDsxhpIqFClAwvWcUGz2WTYIjv5lruOLBIvG0e2FJYJT0MuAr1
Vbb4YSVEZ9eJETPzXLVhFheFrygmIJj38eVc6+/J4nCD6ujsWV/e7PjPuRr7F2mdMI/9JKT1gNsc
5hVjgEyITgpHaC6NeS7E+dUKUHa2LWoUok7LqmJ228e6l3/3nHR37blfal7Ynk7CtCV7ocMoPZIV
zTqi/jhiajDRWXRgAD6V7dXDw4Xc/QB+lENS9Sw0kUEVle4XjX3ZbgHXbxc4H3s+HuxbSzpasbia
YckCytBeUNcatfk48q3X7ktCAzwCn5YWp38fdvCW4y3VEk7eFHuc2CP9gNr5ra6fVq43+dQwGwcc
F5/451aC4omRQlQ90L6G2FKg6eEBwFOu5ZNBJI2so8cEuUGEJ5TIpCDvModO5qp5QKTtSdcasCHK
UBejkNTvP9QiR4DU/As/e7XPXuC+ktoPLNmIXCqe3TRA9phVtvwbE1K3OkI8a+dY4RdbYxL09FYL
KuQ+tVB75aImYbhrJWK7Rtsd2BDuA4hCiLxmdjFRvBAUxDY02A0fi7rsL4EnSLilqEvf+UsF1w+u
RWdV8BMhWtk9BJqNiTfTp76jfLpO9YPiteWZySU3pYNyq3uheqSTAKsyXSiVRFFJLYrpc5vO6X4X
IpedHhdQM0FQR55pe4YcdPeA5SHOmCpL0Sluqtm3pY3ekja+yKzY8vuImfO9shnJnOnZJ2USjkoG
ojIFZVftsnGJVG+C5Wqi8eW+YPzzNjXfeqwStrRvp269zHTGAxSRLNs1Z5X1tVgMbHLVRU8sxfTy
sK7ScLJxqwanC/HNZdWlcMU6C5zaLk8dD5V+ofQC/fggYQW8pFARMEkUjUFyTnrXgVGAgDZCwjJF
rpr+YC01cEW6/XKj6WIiFGPL6o1bDU0uP89bLSDeEJkf+tkvLvV1rQnmdEdz/S/MVRwj3+Pre30O
PhEAUE6a2BQ0keCZUBwLgfmT3k9+fSfYj8+kWUioC0TjP4H+5bmN57gxA8J7PmyiHR1sdGwatqEh
qlp4ZKUPLg+dPiAhHJVFPm44/+qOR4UI9Y9OYyEqNtaVgyIvqE9qy7UILuebpq5/Xf20smUIM7xf
NpulM9e7HOWzYpxwOty5TtUop/PB2184rFwcAt+cozbdf+cFHQjZMhlQ6v8N2vbBvBdPc7hLTygG
9pn7fcXCR00Oxn0Xeb9aQnkc4Ll4HYFTO71l5zz+AgARqvzBqmAgTmjs/a3tBNhT1YLn+KWyj6Ea
dBkPNk6KmxLLjCzg2XP3CyqkAgk4nAUacCse/xUJpbWrmbIvzOVqtxIKHxeSndWwt8KMU5tw0F1P
aUkh0pWJ3n79+mgxHF/IWEVpl+HfEJdVtVIumgV6NXEbjbMBhC2SrY/ntoh14rK4c47Pgl3ff+5W
aAXhHWSgb8Q4x6VCp5AgdhfVjTzsvkcujAvVjzUdkgsTItdu45fFpLIkbbUdQo3bnsybZeJx+gkv
Vc087NUlH9rvKicwnxRCOvUBzlY6uQ9UAl29nwB5Y85tE3NFyQ78tLc6gN5CMMd+R2dvF2xq32B6
5t4EXQ7xmTWg2qFpQnMcX4K2UNSX22Bskx8kYINPbpkrqFGcBcy1GHg4WzutnDcH4Idut8TqEUHj
rE9YQvRa+5uK6ZI1O8Wj1vKT41Cy7h2ceZgLROtHWrskEElGwH/fzSFvMsfrf7AOJ8hvgeH5dBpA
FW0TYFNXdBrOOXcchdBjHcMEjm6XWMqcEvN153IgZA4m6ZZgRQdAHhoOf6JOhQ0aKjHCHYoixANW
sICT8Hor8NPUCLxOSO+0dV06pQmkJUriGS2V/kuRNdomtfT9IpQdLYiOopjc9iM+X9wolK1zPZwC
1opY+A7RxhiAdg0DW5J4E2IpJa7vMMPIkubkbHPYKM5GYSKn4F7u97lsGe21IIN+GFzHWILKrkiN
IO4mFGooDtq4xBoQm2X9P6coeqML7PKPzGWjbKdiqA3LvGOG07dQOcSLHXQ9EGKYCA38zqQuHYZB
6TCqIn0loOm4/+AuiwdgqAZKLwFio+8S3fOSj9GWWOvxW7C5iZnxpj93XQgVC7cYTsyW9cUV5xRZ
9xTW/Hm544xCgJHKFqiJDSEsMAHDUR3nHwtl3LaiI1SN6TaSzKHTqlzIE7VHhutUiRBWIKy/7gAN
jNVGi+d/RXw/FmTGkDhDSItPkJA76zVXhYkwyQOy6+ML5ocRWjtd7N2HCHKe14yIIDGFzDTN+GJJ
bSROzBRPvN7rDY+NaPG7B8mGuE4FL3V3+9uMrwwg7MQvbZOi6clvqAAXrMADxZ+Oq/gY+OFTb6NL
3oLHlvqrzyjNxLrqFQSvFbciw1RYYNqINtSYVmgKm1uAPuC5249N9wLi8WhB0a3f2tZ/8r5g6UhQ
IuSr+PgQ1mP4EO95LGSoBsxf84CzDog5Sn1GdoyvXTCJW9x4edGnfQh0w8GsFJvbfwNi3dh0As2E
MdJ2BRMTfLGJ87v+qYDTFuHA0SLTXJy2WBVCLw9Zhz7EyBFzaFYS6YJ6sytvQvBgQ/Fttj0W8/Ug
nXzbVXVjsglg/SAygZVitD7gmw3fju3jUtSM6F5hAxfP7ZiJPTSWTkNqXzMcRKIWHEl3FCbA+6nh
+EJppBVcKfAhcRg6OLxZCx0SlPyGsrYDAhl1E2DuPHrKXEZRO6XzXScEQKpm2ebuJRAoMmuW2RJS
/Soi3PvUuQY7duswY9P47iIl1V4AgnPjLUpQrdjOOFR3pBsXn/AGuOC+d3+9Rvoi2kok3A9WVnv8
pWfeUYgjFFiGr+ze2fIz78EJrJYM5ehr5lsjswGdlecdvkMnpyF52mY7lKBztdDq4R7+QapLZACm
duYjfEUy6AnvQzmVjdR06fufC4HfUARQoiCsi5yYtbG6NVUTPsl6+pua802i7SPUYpA87z2FfsDn
2cr1TY1Y+3NBrvtZc7Arkp9xPRUaNQ2UrJuvHMFWXx46EQOISPyvm3B7x1gVAAJkUhn9mKEyFPiY
T6l/Ys4LohLLSWX8ttype16FdP/SVLCqLlmdHPeqCI4Gh1F66qVJhRAKpEhgWv7LA42jfcpe7zgi
FJhXs6GKCoHM0abpn/1I9Z2Ghi3d0S7r2PBJftnozTRiNnDWbFsFdi99cCdMMvptw9u8nPoDLPYl
723uO8HkoyKggZxerxXTPWyfc9uE5c6H4jn3hkESBnHuwTsOr2qWgeYQBSSPx76YYP/MCAu3bjj9
cMD+MZjAuF0c2i3skQjr3WacL7ieJcmnl2Q8YbxKsImpjsddXhD43ZgqT/+1XEF577CYn9O2O6kH
B1iiEsavuCXVD0TgKy97OcrQlleUSgSwDTjonEc8kEijIqVsz/IWVacxEnk040/5wIh2vCyXCe2l
yNIC1uCTvnNqb7UTb3+/3Ldp5FLj2OpvuP5s0jMEwDgZyi8Cae5SLkUE+cMzNkr5F43Mzo8IYxJT
nmbojq9sfve4tm9gXF5oKLhVJEiYCvfm134GU/TxRimvctavvzf5YAh7dBq93KcSnprYXchF9mId
AowhKR5WCxrV5rAY+wN/UEgQiINo/3VvmCcAwvjsxlZFZOkVYRwAax5T7b4wnOA5/ix5wXMDleEU
0tofTiUw8ArueFsjyCJTEnaBJelYDW/GP9cJ168+uq528QCHyo4T2oFA8U9UbC98La46LK8ZFCGP
b0tlN6s85iOD/ZosBsICVdXK4vxOOmbgYtbpMEKiVUcHt4MQ6yWvSYBgCyBr3YU1XPDLbm+1CV/g
Jy5t+P0VLt2rIcaAS5jro39TzqnZUkM9HCFguByBnUoJf151qC0JDWAEmEtSI2nnfE2Y5S2p7BFj
fOtTjGMe8gOAb5TzDMdWk1wM5qlFyS3EF1k8a76ksDCmMDaJla0CX9yinUZGKerbE8AcBi+zEijb
OFPlmL5o2gYSVZ2fclCPHZfJRk5bSZkmQTVy0zLP9v6nATxiAIRZ7gcUb7wrWuYmBGbQoxnnEHdc
rcBoQ9WLzTVlxwO7PU26uTCgATNjun1EZ7HZoSr95rINLN2OE7cjcnqzuTkrmVwxppeFNpNJAnBB
JewdyCj1IM8xk0qc2pC7JJB49VrjWxJlkavuLP3JtL8au1bc+dDkyAVCpzj15CCQmdxl8FPMXQD4
MDntMrk7IfuT+7hclPOY2QyfiTxMYJo7VANHSdH4Xr+QysR20ZWD8EWJ+KJcKuQz5JLK3+B73y2L
Ux/HD4h1MB7SYMTd0YtSAdBXDSW6S5PWT0M1nhRPwVCJK1h+0pQ6IwNzqGmZcsc8WLekgJ4HyJrY
BvhIWMbukTWaY62ldtrwlMrs/Dzg1szwYieS6xn8GGgR8Tgk9+SHQX/I5aYVwxkqW3tYTAi7Mg83
P2JQqEM5iRkD2yvrFbLsuWyJfjbsmEQGSQ4FgHs9gD1CuiWt3pFJTJe6syoBUh20dTfvI0MeLNn3
GvmrCExdjuPL7Kmq0ETzCa5cyODayJ8mykpRkJjsI3DwPbjEy/hsvUkZgIuHhdvilzqRNfHrEpGK
eREFDYdjz1lCxgkt3PDs+TK4QnBS5VHvG7aKs46ZY8RDn8ksYTKFg+dEhPm+chilw82A8QKjSnCy
fsfNtyw/HqnAx6yMJindgP0XLEqdigphysbcfUMI4kGMZ/F16zwCjjwL93uP+EKCKWjivhnLWS/v
PZ+ACuUbKT5zPIwSD2o1M1OrLeq379v3wTadCRbm5k42N3XJ81HmeIivOiupaOIYF6fn+YDPu7q0
KqZ9Gh71PrzhM5TouQAi+bHpGDZQjxLIFDgOm+FAlCQ5Irzq6oRmQ2JxXLgzPSHlOIMEQpz92OEL
P+F2JFxlGwf2POjZTE50H+z1uODsB/5Tyd8cc+9oekCc/Gbm84eml0D08wzkn2ULp291z7ByYiLD
xd5qGeFezNvjMwKkLNgj0pQgveci2d23jAnufjsJai1wvYE6eHblQCaFa0NswHcL+C2vB1JGPw+2
M+rWyNEys+hkfFIip1TP0QxGH1jzNWneOiIGT9Q2+J2n7P58x6axa4GWmxcRV1fqrI63F6w9UhIJ
vfmTItcATW33wWn/npCz0L3dbxCFvCOD2cqXJovs/+tMhJ+phVGgX9yCOeOF7H6QIomirVsDdIyP
FjTXdwzte8g5HzqGotIjUPmgN914I0KefYc+I3khSWuZA6HeUkIpUd/E6PnE5aabW8Xchte46gEy
AAFnxVhq4DMK/UPZIRSg1JnZM/S11SRYUnTrdlI8K5WpKh1PSfEkcqdrrWFRWrth8fo1IeSCKnam
jieRF2YmMCWjnfigikw7O2iBFsvgoaPZtOkCmxgiG+EoO6XvonGWvoHtA/co/N5UrLIhsTQ+5R5a
kn/AW0BpSJgZKlvf2B+Uep4i89NJI6FR0guNbvcbDqA3qhuDZFd3Z+DcNva6Q/1Aq9Nha3MZFNbc
4cpE4uTze/aTVdcQ5/O7R9PjcslooPSXr/+F4axKuacHbsGIzJj2lRnJqO2yHnFTvNnu6miNLp10
wiDjrKM1dASomftGbQxp9/MrIpNQIDGxuafEkHl73xMIvCymbYTt9LGmTPIKP7Qb+Vbv+0MZ8lYm
KQQSRPBsTp9VfBxLCkudkinfMxX5Ldhp5v/cYzuGk8JkY04f8NwJW7hhmZ4hh4Wje5vuCu8O5Izu
RcauG/Fnkwd+Qi88FeAWzTkb+1BDyPksMPtYW2szqtrtNuYI1U9GlIkQmvTkfmceFv7tpfpe9ruQ
koQggp9w61tqBGa0QAQ9avOOGs7OKLVVPJZebU5087ukli3cNuQ9dBPMnE47ikBX/5pZ77faoRp+
/uqzHDgy7NueHp01FI/Rx0pvIz5DzlNDQvUbTc2GY1pphlT7RhAsAoganEpwsluYXuM6L3lsT3Bo
s5OMAUP8uX579gqgopcjTp62xsOFK7ZDqwqOwoQGmQ/Hr/9dFOIygtTG5RhhQOHJ3wZPJSV4djnq
03Yy1ABn7z2ny0CLI7hbTA//wDuBrt6Y/3qwtXSBIYEoBpxlFYodCaw9Zmm1qRz6iETLuJJFkonM
/HDCChXvMV8blxwquHAgsRi5l3zRkW38Dm74bZrlVnQRYrvx2cM75/sPl0o/HSBfrPyIoKLIs8B6
hE5Ch9Nz5eaimhEGWIwnNrvNr8cAXT785qgC0EvbsYK8lwTVmYhxJXNBs0KEQGn3bPhVvVEt/4w4
VpYyyljEr9kXMLEJ83YNCAiajtHdCFa/q2fOTG581kAe57VB/ZOEEa7XzYRZdV6vIqCCQNluvjxr
izSvZUJAb+ZUlHkddvyzElHFCjJuDbEDtT0GukmQNLx4Vq5Ha0KzqaQx3wRJUbmlFDXFDLLgZKNe
lTL4z42BbWgPe69meJuKQcOBo7r+vR6exFxroCC+Gf2aCnz5IWlv9+fTiEvo305JktV4nI0V3zkQ
sdn2QTkmhDy4KG87Z1+jMYNC33+cxOMgCagm6QfhxxqZM44SUCn4J95sas4gBPqgJOgQffeBvm4s
kUSndaXjL+VA+e0wD67mUgsOPJEk5VYFOjiufeO8DdoFddftrCsJ9HwG3ljQkQZsbWPuX6KjipVr
Gd2fcSQM2+WTvAfLEJ3iLoz4Ob1ToUr6L4WpQ0tus0PJH+aTlPzmo52tM31o6mYaMhsVrgbJ7OOm
orSSJ9dIsZwVmXdCtxnq+9xNVCGCJd3mcjJWm3qOQkmdtXaQeaThsqjYCDEaBzVg8FKvecwiBVEb
LFET3mJ8uAdeGcwOMmqDxTtl1sYnFySHN3VNS8eEyZifb7UvjYsPn752mLvN0PO5jUDkmSMlIPEJ
DzQYfeypViGASCg6v5QkwMW/1gi8il7IRDBW9xKAQmZxcje/hA+5wQDTQAJZfvErMMypddG82LuG
0C2dN977vCNYyWhujTvhmew8wkztDbww3sL03/hiPNANDjJPZ8bkBjdj4ADJ13kWi3gZtf+Ni6i5
o2gc09DLn4ejccfp2+e76dZOOxH/4lBMj90I60tLXbqnr4W7PXJpzL1UHURRy0SssD+cGheTGRzj
AJ4Ss1h1jRKfENyW22GoZ4ne8QhzBxoAwVdXz4WPgNolypYWLzrsepcoxwlhhVgkxO/ijx3cRuMB
hNpv92w0m+MSuirDIWeV0zwsR60jHwKIMmBveVS0KPZMO/lci19LZ2355BctSmOrvHZz75IA+KpH
bs5BSgwHX43QKMr35pFxaCfNDUYOLz2jeCaMFe8tI+CM5jji0D0wKLAGGs7bsduVw1JSSbzfHHMi
1qIuRtEWCbGrWtuwbBDTYztfYQeEf5uaHtEl8aRxx1d36//ruK3vMymkXmcQeB77FllZWSgJ9Psd
VMrE3KNZC+e1Jw7uFW02zZiI8WmrCNEkSBsgMPftfakaSXrVTNpRdAyaWn80jrT8EavhAx7lgGhs
Vca/ty7tvvt0yE8NYOrZxXf6/AbOsYoVv6QOGdyeTT5zT1vBPD1c2akWKiVUaLuVcQBMFI+ArgCq
kGMIZUpb/+NsPibjM6WpKIg0ZvPhaFd3BAXiGuj/q2/T7J2ZKzCapdrqa1Bzo1KW/FYiiJZ+sm+A
iciYc+HJr7FmkIvkcduYxqK/SkmRBO8K+f9KHvkwl/jolLhw7Pc8nciGsFvZdEjZWgrIHAF6lNuK
GRD0a+RTK4YZKnPQHRQuYBho6cC+VqckIqUpz5rI/2NjQ+53JkqVW1tECQ4Qx0+HPG5IbOSSngQw
ksNwv/SyoheW4n8Rb0nElOdOIniDLtCdq7UWgJMdSrt39Ja3x0nS+VceHXcnEVvZ9qjuaFOWtVUw
BPllRjQ8XgVDIHmGDDAsAYE47z2IXNDzoJ6T+07dYbBSFrK01QnHiPtNTSQYgpLtkeziXseB8m/e
K26G5CZNAAtn8R5TCFOg6jv49LKHBZa97ZmaYAqOmS3WRP/7CNHNItLGpIFGZFC6J4gUHXJQw4HT
QbSwVhYkhbquqOnOrTjl/UrNfrgSeqkncv2criOLszjhiCfrLdhwgtELBdywGDO/ivWvuuX6R1vO
pro4hCiO4siVYk4xCqC7kmzUMwkb1FP3BW3lQMYeMHcPrF/PXWF3/lcE1StQ7xiSEbKf1gXszBQC
2cX79gJhmYslDBuIW/1FQXV1tDc4PLD1lD9rOyQcgnYeGRCrEHlXd4WnNnotqLddgHrIyuEbCLoh
VJqqla2D3mf2j6hp8kkKWtnKEuBJw/axbToDJLPJ8qt2IaYRoY3ZX87WEFx403e5GtTLAGwTHzYX
FxER14a4gKzK79KlkOr0HDqMzP1AVTsFtYKMd818ImiMKVsFzXfe9Zf5vg1jNFQw4RVoOyKx2Pgn
AV4RgIJe16KeA3r/qJvaju0u2Nn5yaFh+WWGy9x+1oiPkE+/4XTLk9kuaPkBK8ns+NWFRdZ6ySCg
YmTT4kg0pFxUASj2ED1C+YEJOugIrE7q8CCoDE80xjxS4FPiTyc/6zJ6tZ9mqdbaLQuboaGCHAJ/
t1lddARuug02CY1sTJGTaumMylur0/ZK48REIbR4uabnDd780zpR49jyhYt6UctFH7gneBPzoNsh
FkxX9ErvZuiGCI2iIAByGHASOgcaqb4U4TEmf6ts2sOghHTnfEG8ZVULf2NFKgWoFRP2OCWzd93W
PW3D0RAMtsE+98DsQKz90ushVGVTJmV67T+v4zpnwe2UmxGQeYgn43qlcG39JU+UlTNxE6QXCJ/w
+xRDZTpO7nyxxa77NhDED00fEoET1Wg3/fg48mOHCTmbfnHoBj9i8z5QpPoE/Xig6p1V+2RHbiiv
xot6wS+6LBlZGGHTMNSccS8mZhBYie2WRL5ZmHF+O2O2DjKoETOKu+By8rhhmoZbj12HyOYBuHnC
hqGpnDJUbnhP1VQA2NEypCdWElpxv+ya/2R9k8cfBohYFZewi4afL6Z13+0EWT/OnBwOOq5wj+Nz
w32mXq2lMfCjoCVCfPYs8Q3j2ueAbGba05cZ4fIs8+Dm8/J/0bHDfEdunRE50P4feBdNIA6PFQAS
b1imn3Dibiujp3fw4n9D4EfE1kd8ufUQTuWxrJoMoUCLiFRwCSnQjrdNi6730V3+/FLSdsqmlFKU
4ImjEbctzgwHxNi7lX+EsgAbvHlGPiN1cY6JfF6Q9dgWNBQAlWLXE5NfWMAIaIeezNxUucehtuiA
t4e41PhaBSqcWGVpQQuMx4g8g1W5a/dOn/XdXyzs/MuZ1fHVFtxaY3ovgIc+fTRUnu02spReFtcj
aKaS84F/krKHtTHXvAC4oVDKxJAnCV4N8dowh5cceJznfXjT5Fysj3BAitgNNB7Kb3xUkRtJ5TKk
qI+ahCZVUkj/Uz7d/kKqcHbb8tiq6BvhC8ZhVhb4exeXKOmZ4jM6r+dPJskWuaPAgg6bIR4f4RuA
KCMOeQvRIHfuI5CGUorn2A6lnuRytJp7PY2xisoqik7vKSkGixbEajdPbDA1o4oCw54pTpG/IHMf
TymItfPVCqSHdrvZAjdvzv1GVkBFYfc5Fk73dXSRe308gpnFqBlSoyKyuGrnopzqdTov78DWB7iz
ZAk0uqzhCaH52U3Rb1lsPjchTk8SX/OWL+pmM746efBi42qNWComcBdrSQ3zmTj2BGVpVg6loVF3
cP9B5baZOGsh4qLsx1ZZss0M/6jiOfXWLBe6ICLZH8eBvbnQfSjJsm41qJ1yzwdFHcMFuGX1M2OZ
DoWMK5t8pGOg0Lypw3RXnydCvxclBbnobpKzIL/xFtAuVc9ibledrhFXwEcSiQH8cOtUFv6cz7ag
MbDLRve7Z+bUhCw5li5BgeEN7uEA2gCAq08gSv4XJWZ7NxBRY4CQOYreRUTmxKSXcFSAWeA7hBtL
8W0P38vM/KZvPB9IhZ6npTW8XNVK6e6CWO/AOMjLHm0wYn8huBax7Hpc7quP1YxogrQsr3ybYntk
OfABpzBgMDNLlsOnmlx8q+ybOpmZM5+9LiSShOtudxdWG5BxWd1Fl79JhzREkFJ4Y+rx8rfQPwse
g5XYt6IrqRYUqKeFsf1hO2QEKgIk5tJFJj8GcLrRzK+LLHmeXGgFVkyGH/BfwS5lBf3ZO744C0/D
GJ3nbyti8P47i+HUla+62wBZ4BNtG00kEpr5Qesu7ACIn/9mzIE7NBiW++zHb1+7Bk+0zvssidLz
fssf2I3uSwnl+fp6csEQxKZLOGezhaEMBpHJiceEVWNlGj53p9k7HbMFnPWhvabnoXcsj7lFJBBy
78a5JuqbFLVIjW2Mh8BwgeMArQ0sGFoyKGl/bKJyqwBWzqZ3NOkid7H7X6JRJT5qE3+ezht1Z0G2
2u9lQ+GR2/IQq3C8yHTFg3h5X1iZic5ARIHgPD9MZ3Yz1Z9cZCjQdNF8czikh47uJqkK2yTBXxlH
EzZvCjiBFv6nxc0QbfJlX3vlsiShU9APGBcrW8NN1yYKSRaFwdYoLn/0TmmGnCBYvYdQl0TLvBV7
xqTvRIqWeT9VOgWw/gM9AxzwFnBlwS0tOAGIdv/cm6vUKqzQGMNj0Rx5/wDzE4iI4uew5wca/f9u
DtNQ4+/NR2RnVgSMxROkA4+ZphtMQhTuuo17QFxKkOcSPA6MoDRZDjlLPY2ue5F3n9QFpuZxfBIJ
iLDtWAmrDA6s55XhWThBz0eoFaQ4u9Jatcm5s5W/x95v6bCJ/oOR8A2frKuE/TJLNinXkKX96vNz
sbgi+ezgLYxGl/QwWu4lN/j1fHm4Cvl+oTRx17pVYpHzS/6WsberXm1YZiFCjA7TLrvJf8DuwMi4
HJ7hrBqHp5SguM1PJJiQ8DfmMjUsus/enXYOzP6QrxZBboZ7F1S0AoqjsDA9Y74j46IfcnXRkjVX
Jfk3OgS5+c6Ph/XFH+VS377BrshdKOOPuvENsf7kV9cKmkWwFwcXMdtxWP6XdiWD0cW9JN1hDfOR
MZDCm8cKIfSnrWW5vRRkrNwRTcE5v+kCAs7pGI8EanMx2tof7cOUZo2zIPUvzqyLCw9vk6qpKPof
qxv0+NZk3aHLFaYeEt/faw2N5yBYcyjoU/Gl2vj7sib6lnagnI+IXffbgnqmGpGa5uuZJ+J4qLWJ
3n3dB4H4wbrEeGXGXEGGLBO90l4fffTbkYXVz766b9SVdIz+3hlSuh5UITddkvFzRACRviM/e1qb
aMkeIKnHw1OGYiP0enyeScQ5nir+vO2WbuJw27MsDkSWfWCnfuGFV02wIArWOZPcbcVATtTDL1S5
yRvsM7g2s6UeSfnG5aa18QWLo2NN5XuK2yRl1/7tTUjDBmBoXLZEd6Byt3T9aQoT8wRgaiMn8wpV
oQiRR4jEz3B624sGALZIWhEMzGd3SIkqg5EL/LW5WNK5tyAI+rD9my30TN4IiW224dv1niO1qM5E
hkC1l/YW7PO8IKT4JGGA5EOZ2aEQUXvAwiU4bYXdd+Pw24RR2tNA3skpjRBBypZEcMOo6b6VDtSP
vKjst3FMZTfgwnvb1vJWqonCusD+/ehqrBi9q9FijvAVR7nC7iWcy5TxCuKC0GCoWcoIJU33LVe4
J8cDoAdyqbRttXWMlHpBtbsuRU+QTNeypcETbSNwYtP2HCZ/fxfmyblyw8WuDf1jRyUisGX71Ckn
qJjWrX0VKv5zi6eAc8qqHE0RNQOWBzBQS1GW9378PQYYBFSO0klXNg/F6M3fznItVtnkh0IDhDzk
M9C8hfuYRvrP0H9GIHLNuhjYE/Q6k2A0B7elOd117V3FmDpcSwYTIfx18Mg2dtKYZgEoLlojPQ4O
3pdknzXnYXvWEnP/oU+oLy2T/xC+0sPI1kWwhOgNfPet0kpakrqSq84X7tpdVKzr1y6oHhIcQfBM
gBfO7uDtmZKeWFzt0+3F2s/tLZ9CCdC6S2fSjIR8jVbvXz8bpevnehBtjMx9zoYuQ8YIOaanElyU
8xH532onIeDlh9Cun2uK1JDw8F7/bMebpjGzxmupX2s+8evb7UO5E+fqZZ7aV5G6iYHvoPJTYa0T
I8Or+u/A4+wPrs+KfWbdpq3mUFpIwoB08vg7//rKc8kYXrF/LC8WmFFCtH8/q+i7INZYbYvZPv6D
PbfvLkobBUPb57Hcy24xuMzmKUzDkcVXoXQsT8jrHoquQoacVzIfpWuTsubAQM57jMY/sjKBAPvp
ZNBZNQr80uhpZWc8BNv12X/ijDYMbqVrNf5ZKdmkHFOEcye6eE3HWzdEnwts3d7uza9TClrEgewm
pHdaXRX/WmgUjr81oXhQ31TKg1JXyKfwhKOy6iDT2zhxXS7StA4KR32bUEg3q4mXQjwM3/BD1Msh
+4JSk/7E9Odil9Y2i/tYnkV2j85Fl9mTqvdpBGmTkTKTnEnztdjDzUlqJBXHZ6mgFBr/ryNZUXiP
d1nRhtwYvA9Rdl3cdQPsuKa6RAlbHMX39QpkQ3x6hA6QPbu6h9KyX1KK/U8DfQhv9wlQ5Of0SDll
x/bdJsyW8il28v6wttETOGPp+N9m08K3YXU1jaYSexOuyH2nzMFIZZLx47uS6O+ql38nOMN4fdKx
DfgNv4ZJHj2QWBzzdJ444m40u7mqAUKEiw+JFHKASH3I7tqamMohtpYiTzjr5RzFNHDdozVmFCTp
neWP8iWVYcjpuYFropp98SE46I0scRike06lGEiqiSZiKzPNK4u5EUmkSi//HwqkCZbTJvaQ4QMv
PWUya2AqW1SFC4uJ5fO84o5XWDG4QWdokLtihqSALehUbZtJu/kw3fZ+mjziw5aIfCqJXXLDYEPT
VgRp7bStuLrD6rnPiLYpi6l3RFKa17rqQadcxdls9p3hp7aNCLiE9pPWYXBCQF3t/bOKiIZpRAmS
fXvj/y3HhBtu67SV/hi0hoIj+GHQiFME2pS9fWE4FsbcMf/nZDEAMK4RQllFQuolb2TvJDK9ME8M
T2PSvcMPBUkyUt4YbIh9oGx4CZi55aYcoT2tRnEiXJ3I3OIZQHx5W5Sz/y4XhwJeZmkjaNrj5WL4
rq+w14deby5wzPiJUBK7r6OEzt8w/ZfKXTt4FV7XK8BpXS4YUI5d0xf1Ok1psTF+0RWb04E7zyXd
kvNLhbwLoOcYbLJrwDZjhvx5OjYuyK3KxikCLB454ww1WXS4q0GcO8A4WTFH9uX6Hk4IwBsPuLcn
sXF4QfCNbHWkalYanaHtTvVFOWF9OYU0ZS0JyRbPyrX11ArWbPB5Oro11gzIyC4AoTr9Inby3Wag
e9EP6pHocfvXp5rx94FKxvc2eYcReCufJLfFzMDeZod9+DHXFQ+1rIaJA10NhNKIZGIXi+5Pp1tC
9TQeq2N6teRQ5iHIlP0DjWyc6ordrZe5npxNjbtttzWwJN6QQ8sEfgD7aVvA+5QEDrSsNncS977K
KO1Fbv6EQZQOoB6AsA77F/tT16xuyMWjlmqHkgU6Z0zXwcJO+AQMgDDjctjTJnwjrE9bicJcVlgK
dh+Rgb9Ozs7/Pp+kBk81Lx2kaP6Nzy22cDLmPHjDz+R7ZJtTXA0zuSwI847gjVcFmpHUy9/VQwxV
iRV21tR6KW7lTKnvm3DyWNRStExSNlluTJ86RmnD/edynLm/nJzOeWC0MLmTQ90JkmZcffraIVxh
3e5uC4dkE6OUw8A88TUhQZRN/GtckbsrFu8xQWJn/GmNsV7bWN5af0Sm7NZnoiRabrky9dCmZ5XM
0yV9uDspCIl85iAcDziLAubkdUw2KG+lPkdU3/ctwDakIlJZfdIJ+BRoy+8RlrFRJtXDlzRP7YJu
fMf7+traMoCTzR5pYIxza8mwxuuZTqxT1E8JHKWp0hcgHPvYvULvlMu4P0mXVEvAKZ17ucndysf3
QFp4eEn+pDGWIuCxjYDfdbYR9iDyL3jMphQt1NkaJEFXoh/jA5/9eDXE91L6HZKNYWtwfmHs/YyN
UT4Xt2SLH4We0hq1h0f0Hxf5sxfj0eqvJ48xeXTqXdI2Y6rMSkCPXkVRO8s7jm5OiUUd1qThhuPj
+l3RnVUCfBfiP65/dG2iGi0/TJ0cbCGZn6w88ayUh3naWG/2QtGcnbDLCWYczIkBne3KNfsg04vB
KaUDOBj61re6pAcDeE2Ygr70ZaBlkxPijRgl3eTDyisD6wmRJWgdIyGCR16tnCdIT9TG2h+pKHw7
Q9LzH4uDyPnMuG+Q6LopBGdN4MCnH4cVHCEMZ1q2Wd0s0sHFLV2QLT3k/G+Y9BRwJjeoDL+BBebh
RaMISq53d1dCsW7jnDh5tRkk4ie0IsxszWaTsjzJY2s4hS2JoADao1RQrzM6f0sOCUXOMSv//+j1
yXbaZnhMe9k7brRn5ntg61lKpBAhiNUTwq404lSfV5kWjIJk6wi3z7gB5jpGaSUE9QAMj0ENnI9Y
d4QULUSUQLEj4+vr1NVUei9B4zeD0/crLEhFO6Ho+QvoOIRpmsBuBYFu52vuAs2eqL1cQBxD66uX
EPTVH0gODNk7CZ7+HK98LFB8XvQTziSt+puROFXGlboUj5af+oj1fASH+UAsIYh4/RyeKNo0Cah+
Mw9atHCBzVDTwCY9oGbXKuJop1qHLW1gwmYXAa7hl2YT7PFVtfrlk3JGPZCjam/X6wXS89CQKGFn
ahK+a1j8tyIAHXbjqTaf2SNMP9LQAKaUUVp7nBET7v/5RFOzcp4AD7nWD+qtDTAeTngEsHQUBg1G
jJ2GzmAtNRoF3dCv2RSFpSmHQ6qI8u1qKorqvdjjlyGMTxyqO4Z5eFWpRAmVAiGVu7CGnNtVa0lo
pm3AnvPl0K/3UDzuFNUy5s1F9RKpHL3ekTJXn/Hr5+qICHeuROqMuw06w0KNrc+jSIu/zV6VY1fr
cCxN37s7kB/tqo4qCmTkU3+n4SKK9ull4sT2r7juH6cLx2CT+1ap9MGeLgrDp/sqkmc6KYe8yOkD
KjEMw5G2HOdt0ODQw9zYc9iIrI03BWsNUH/BvV/ZQIgnI9P/Lli5BPZT9K8j0iaGCgypqnQTYEik
CKVZ7a+66YMvgfdzeSSJany66nG8jk/6iW3E9sxygCmvjSBFwcP1AyGSc+7UU9Oy/WAX7UpxuOC3
wu6b5voz7UwRu/xvXKlWuDEJYfjipxDE907rJTH8GAsPzkos7ehN9xLkZEmgepYZSo5AqTz4Khmc
aKG5/4w3Zt0q25g1UVaewGqMSxhwJLyESQMN/MPDaRIYM2sYtJw/x3+Yw3YcORs42dyqtyfE9qqG
TxolD/y6Ll8Z4Xp8jXLhjGjyx0uS01NkkZI2UjuGJau70oxzHxY2Z+bkkQsNkjDe7fSioCITD8JL
Ym7p08sftG5smMOswSVQDZuzO5+RGKEbc2IzFDLdlwDqe/KT40GGpjqwEHyRAQ4SWIkL/hvIZqSU
SrKyf1XML3cGpzAbPnh91LhM34AXfU1PNfY7zeBQa7qdyrlBqwFmyCTl1HHdYCd1gDYpD0MzoLbL
CGhkhWuVfxEuo7BUQ3Lw2/Bl51GumDt27oxfa9qm1GFXAvwTUxHALJnMha96BYTlq569bYSDR+nv
9lR3zARluS1g9P7xbF77ZFpWb/rvGDbWy1C8Q1I1VQEAICYAZ7sM+weEkWFD5Mta2MvhNkZZKYA3
eoy2laAvfjdqjJmdtb59IArTUPFG7fS5E3MLk0D+rFzVncJ7DG+5SbZ5+sDFj+NPvthM8pHbRs6e
VK3/M3DeGaEySRMhMkrAJ1IqlxIJpsdahFC9WbMTN6iLXGX0dK6A6mLnNqXEUQ0leaLtuzyJZ02U
8Gp72DnBDJnu3YWu8NKg+shiKPnjYzBmRcK/V5XRuo05QePa+1Ta4HEuq6SbLSdR/QUpmJOdGnWs
/x/wLPlgSYVUtalSYHjVjXPY1a5HZ/yaFOvFk6QQg0/QCulfXpj0wDnvUDZ6P/TlsiaUOE3cBP75
1CfbHbDJxV2OkSITZHZpa2ZI2X13zYy2xSZJ+FonpkcCrvbdntf28ZyHB5gVnRqEjpszRKVnpyck
lQzBnXh9fimWhVnTHRoyuyhU5TbQwVEKka+w3qYzIOxHWAO3rAhpXoKe6qNiypg4IqfitMVlkKdo
CWm6CrEx0LH6yZj/BsiFblTnt4QbLyXn3veD6lcRQqBr5C8/0crYgTbwDH/ALGKY1Mo8z34Y9WJF
medkNjmiSeOQDhTkm2K+/HQcH6mRFokxlkAIsERRXl3TuDfrtwk2gUVoLX6QcpP0dlUGG2QjpD69
6CPmhI4qyCmLVe8yKIx6rSa4L1ErUdRnRHH4Gq8eyg5Ffvr5kOhCMtXaxQ234dn/eg0oSkQn8uyw
E71rHGyg8xGpYwEkQ+85edL6xAdmLfCuIOv7o+bE0YQWlrnGpyTa730aL2VzbdCB8FIRxeZzBP1W
T8mLvO1vZIuiAmZTDPPaGLTSUweVy519e1/HQ0SK8YVrBp/hGWkcY/Yq8H53SU4RTPgKlSlK9/xp
rGznd2T6kAuVhaGYYmgcM3N0l4yb+BGkGDaDF8SE++6YuKJ0YKxEB5DISQxkV/97JXURReRedcXc
i7htzLjUdpwEAe+p6xFQRe/imUfn7k9f845QOQsJ2gYVKE1qbSM2Fr/cqIAQaTfwtllgFCCwo7/1
g+ItMoXCwo8xu1D62z2I5xYqUFaJYSGRKbQ6RhQa0zuQO9RjYin6u3GZtHS3YF0MBmw4NDrtWws9
zYMEjfwCnhRhT1aHT+NSS2egOQJfWCeLOM4Li1zjEDhE9w0HGgIfxQ/doLbFRdAkkA7fHh4C2U5z
mWx/I9Q9WeZL8qaPwytLIveH3FbsZEk0Lo4+koULSIJW7lMkscpt4mAAQu3vfPYZu92W9mT6phQc
loXr9dwYc+yzcoBhCU+zdAI9IgwqiYQA/M9xT/JATSTkfJmyRxCheiuDmY/Sjq0vFt4RVb3ZiCtT
mRXgjNuFHgxaZpYtFAizKLeCdnLvPcCBpVsI4ckBbtzlZ0cJp5PHMs0TKEU04UhORcZunPX4L70M
X+1GRsYU3Px10H1Pty4zs9gBtFOGFbslUzJRP1oxRPLPOSnfEDlYDFxe6e+z0t3yVrtWADCRlibr
ReET9E6PcsV/KMcagvHzfO3F/QEypiVfJUof0lMzpYWVYW6ilodDexXbiKUU032jVbAiV53NZyZC
XiwlbOBN8Vpbs1dkfZc97fOKjGCtewHOFCcimE9xgEGXoQvIConJPiNiZV5b/i6iJftDQcyar0OT
qLp3InBNSAYNWpnxdyVMonIKWUw8C6UYcm+78yKFYtSp3Qcb5hlDdHlmObgLCvmI8kkr+f4PHVzS
oxrnv9EmYYAm43HVAkDaoE60RUI2y86O+LdMRF0TJx8RviMp7++wn+6SmXxX26QOpx0C3ujSVO6k
eDJ5US/ReacnHvkg9OPdwcnEEakXmuqMIz9dU4tV1WlmnrH3JPmvp6mM8/dz6PWxRAPu5Fu+3Fu2
WCUcSyGVmwUVnPjH/D5OUJLH61sJb9UzT6OmZyJRLqNxFRBHYWfQl9mhh69S2izvdtFEWTrsCUqa
87XGoGJjfmDmvIRAIXszH1SbYDXLKn8t+HI7SqSlc6Y4/eqtEzC2BqE+7jcB31RBl/bOvO6PIgGL
YqGkG7QSVV0pJzSMt8vBBEnFtHGxXrSi3wZa0n+E1aUoR+idO5CRkXm3e/oBVbev9ik4N6SQHG48
8akaYy+GkYplgps0l5HPSocjBTibZK7ZMjigngdxutS85yUBaV0b3aiw+dT8vJ+CW1Ayzj+Mr4da
JmsdufVvhvSKNwX30y8Mn1p9P0/yeuFJY9JEFAN9XYNWHJNzKkvvufauf+CjnZ3TCRDl7fwwLLOh
D9ozk4h/XV7ACLLkcjHzJOcPKAvYTlzlJ1t589DqwYSgYd/LIaJqQVwQms7bPCFEZKdSZ4tY0zOZ
REV/vVlORQsH4B2cdXfDgmj6Oggo4PSj6jkU0d3ZSTH/S5Cc+N8ThvFAu8eLVsVAs/ElTLKv5bom
HMz7gvSBtiJ+X3DD8fzF3aQDNwE9fi65FGC+CLRCp8v7jNKMgCAbc82EqYoIgO3mMmqWjndL0gtl
RwThTLm+ToDytlu3tzM/QeeXT99oCrvc2LI7LeOHKVMG3CVN3f9AizR+sjn85xzIoELq46g0TCAM
dA2e1bhgO/H9PmAPkbjblAzRDw4jNuix9LNpPXWWlTunDCCnQSDeNyYaGhtlGDSkTb5lC65oOPvj
wUMuRtGoPePADwat/SxaY036zRhwy6i2Q964Dl3CVVRMuRSrnncsfPV5FRH7GC6WAwfmDuirRT6j
VEUzrgAWgz8eT4S/4kiDWWhmgOBZ+ZuxssYXMfDdqvog+yi9kFE1HmeB7vn2TLDixY6CaAUisczN
zsNPYV2nPnV8BWrtzYQyHhFdvWTpKtvcAZ3m31PeLRMx76aTPDOPxmxr5DAlku/x6azx6rhkAdsu
zPrBJ1cPuPt33L3HghSc+fv58BwUQh+RULSCs7IwXx1pY5O/vt0HyArwm5v0h333OmSAnQOnau5b
2fDn283aVhv3+kmr6ddiA50Ow7UDZG4bsoIQbnLLUpEr1xutolxp8/XA7hC64eCMGkTOQ6pJxexF
0gDMSPtmpO+XYwo8AM5gIT+FGrUceaJAf5Dj2b2TrISTWjHKVO5gmpR+QrGjbHE9bdNHwTfPEJTv
Qbqj+Io2vcVWWnYic50vAAPnrjNL7VSQEQNI25Z9bL7ne1STjDteiIXnP9+jTbkkEdHq83XKmcsE
/4nzhoK0lJ+ltIYgV7juhBYQk6kzfQiIlfE/pCuvIsxTiXO6lT/2WlnSTj2L2BAVpWM+yJeYQ8sD
A4QUi5OShb9/eD5qGXYpEbsBJo2j2D1RojjwegHtZrefOYRXXbgClpnDnu7PAX3Czg+1ZjMHug9O
vvAPPjzCmEpETJW6aH3WjeC1W/uxgYDc6rM883ZZWZeU6ZTYzoZ3ddKv7d/j46gtyfkv+C1EiIBc
HSjPJmLF+4WJeIKiMoEqiL2NWUWoyyAvw+VD5QniRdhCh++X52ZA94QyG98zevWjvULqUcI8YEEX
hLPBLrU6k9ZkdEH4M726yo+oQS+ZtZs+wwyZjQN4W6UXxTgxy8zqT8/3QDhp3wVP8PSvo6+AmMUn
LrYvrygoTymeNoS7Twv5kAYiwmp7HWzmi9DGRfNjPpvY9FLXlnoQEKrRDmbR7AUH1AvsZ8dd9Yaw
7j5lNAkt7poLXHlJGrqrI1D0QgcgpWoIct74eE4rC1w0zvhbJm7TnlYj9oG2XXpkjTCrz13Rt7FU
1qPPtfasrNh8zhYjmuS6vYuuOYfaDmOG/5lOoIxt6+H1Up5bUL84t5jXEgR7FJURnxUHkJdkMHdf
s042L2DOaFtkETeQzTeH1TpmPZQHZarLUhXJtAfRhLS4fuh2yt5UkZ7TyXmlbtLkh6QS/x4YHcD5
i2puTUAJJhkygaLmSNsG95XzWSvgFAAfWAJYxkEiNwaDD4SQEjXW8qIFApDOsedRMyYJPgaQuju4
xmaWVaacgDUVu+DvsdZ7VDRHlicO2DMXvAdaq+XQlKGkUDunVkGsE3nBTuBcm3rnJWFMiQi4RnrY
tUaq1/0LSix+nRfQGuMZ9ra2GcmQityv9bgpxbj3gWUWIJvfqY3GxaBQkBPrXPn2buWHY7nZ1Y16
kHCKjNJXpYujkB4FU0riUWsJ8FOJmJjKQMmxcaYJEg+XaB93pYhUe6iQjn9LAmV7ZoGETo3OrV1f
53QmhIMJV3atDfPbCV0Orzay6Ma7N07gwhO9Rxpff4Hop97HCbbHoS3/q6c5bXZIPGTaFWTpcaVk
M+2t90+sbG7QdCkPjM/0B71A8UaI3i0HjBAQBjyvQPjWE43dvCiQtHrvYD3brp7S19ax0DRsbzMh
wDikU/N2a5Y6IE2olIj0kQZmrVpM1Tp41i28ua4VrHj1UCk+vkO9MR0HIo8ohCedCu8hLd19bN60
Fy1jb6xw0aEi5/JW/EGZmHaxoioFHPavIDSEr88N6L2vTxmywbcr8PxcqWR1LY+kzGo4kxJ6vbUW
dT/eZbA+SbLd+Q787pVuQbzVI+Cfxmi9JnnrzelU+XqWbIyaimPiXT+G8ETfvQhEHMSFULNDG2Iq
tOkIisLzg+ciinccTD/eH13acr2Dk4/r48D9z6nTU0J7QAUJJ8vUP0qTlzoK8hB1Idgy1QqVdXna
9n8LKwINzE7vxSo+u/kzPix/97CLZGlhNhrcfGhfUeh+9wBXv6a24wrPFM63q+pP7Z1FD9eQteYN
DndK/SjxuJTpNSpuVPhHv9HoM62R+9DhKVLnn4qpq9y6oALvemiUArrOGAaPSj6RaYvE3ayLvmLe
QGBwtA3SteLZl3yJDUA9vZ3VhME+PMT8EL/3zCIz6U/gvf0fqL4eRpMRAEUf0MnlGpAM3XORZaoS
6hDBAnV5ujPiA7wpsXfGtRoE+2uvP060IxhO99+JZF3ifQGyCSPvJ0ipIF2/HWHFWhY+1ZYcHnqs
t/v0TuVNjf7N2PR+PECvv4+rNbcPjaobDtAnqW2szHA82yY5hVXplF5RpsELdmfVhE6yc1sYN47M
Q7O6xgw0Y4ocVQBe3v2SrPoj6FiIl+fTNScmcZbBxt1STD9AzyBZZsZyoaplOK05YGGWy0eG/2B3
E9wUqd08aDQTcKY/d8VCvkbMzFoVz6iG/lcdreiVBB4s/PJXH3G6dBhOtOdMLt8jNo+aHnIVkcVk
1ZJAl6XaHpg+8JsuN85igKeCeaZ7bUkz9QFqwEWneRJQM0KV9cY8hn9EZ73ixfWuviDYgstf3IMp
ugdM+1E/4xYTdr4ky0iIhD5mQCp7GBSmFFXGpbF0k9C2w0rFPXcdlWQO2FTNA7LMaC/EG3FF9uXk
LZkcSjwy1eLU22nYOQlbPFYivL0px3no6nW9ymrH+WlrZs3Q5epIvG1PnmyEveaG8h5tjlsONzFi
mUcGfEXGBWOlrD9ria5RZiObd37xKHVKLHe9IjhDqSV3a+52st/+1zTZpzFcqoPtTlgUKC1brp1w
JxtswYe03TJHVJsQdjOYZ6oj1Z3T9ty++FoUvckMI3lqnekl8DM2iG9lHXoHJ2o/NVXy6bjH46pZ
3OI4lzZBznjjqSXl8hqo1SAGSztlgGLh4FEEuI8C8DS6Os0kjhsmxfFEwCgWEoz6i5AmZDi9cnNI
tGyW7QspkM7yrSkbZ/Rx0P03fsFzFzPBMgsfcObHJEI385hgh1wDkdM+tXr8hjDVbAQJz+G7Np3K
zUu4Khm+xUCZZY6eYdQW9zLILrAbVZKv71mVSHaTxwHFzs8v36xEoFf/a9vhjrL3ld25ackoJ2A1
clJM5zbwjDNEqC3gE34/tJn2CZMtORAc/6fos6cdEwNF+HYZdclvVd6DPFkKTduCct+MfF/vfhqb
BMeT7IdChvw2VnNsY5bChSo6VpB7RS9xXGescg5WYXmYGk3/9hLfHrVS5zaRe0tiaQXVZiRoe2qg
IzUE/qRdJ2PQ3nYtGRhZlxRhbx56HjjHEieBWkuF+Xa0XEfpvqdAyBDCN1bqGgmAKWM9sepEUSo7
moqCD4+2D1N8VVXgPAvZkWumFhPUJ8VppXNhkNNiuLevdMRwayVsgFqVsL2OPd5aJz52ebwnyQDm
jaavU0xGTJ43GMTkXDHQ+7TMesoaxr4MZKjTgs8EF+e0Wj7gGVpkjzFAWRbjlMn5WHQG/w3Vt2mC
RkSWcNPQaW9SFOjqTaVKsMpzbJGGDfjIPTDykfyxR/+ENPhhYq4pO5QaFQ/DmmFn1uZlxP63AO6+
NoffE5za6e18iRDhlmYM/1X+wjTIqM8dQAhpsSkpDhPGTA7AiGYdlKlYSN/Y9OmhBew2wTp/F4yc
0eC9JubAEt7kLFOpKO4wdH8elOxIzDYhdKlsG1hs7Bnh0iyhOIsIi/KKzMdOHGw2tvpe7E1dqyss
gQYErTavFLlI7Yc8bpJm8E4v8PZXBfRR1qARWJpyyVWpCnPC+2j1q+86KEjbZWphiG7+BLSVvkKb
GQMB34bJxM9UmB1YzTnf5bq1+FovVrdqNhEpjA7IVPrYa+/Z+KowTr0fVkJJxqoAcKIbriNhO+70
r82JzUCPy8U2lONW53naG9hkhXunEnl8SMu2tzVtG7HyA76Y9lhWK6MrA9YLrffl3/c2lVDiDMQI
BL49Q0WaG/56PNVfSEtXDxOw6svKdjURdFt/HVA+yjOUzcCLXbBpFWj65M3AVgBGsrJNKpCnc/am
p/LzHJ+LdPluUxgMFf3xaAXJ5ruCSNpeHLkIT6sa2RXm5l2Vkk1O0zNCQsc7nva8O5fVsF6HAF1Q
W2ow6Xp1iGlMetiStxMy9LKasOhc732M599L+4KKau8z/2zBL0lhuX+kyQf9Ji0Va4UrrKs4R0Zk
awxreM48f26mVrrojOh1VSGV0qnJqfdCssynZVlUZiD4wFh3M1WgaBV4XTGvxjaoicP40bsXiphw
PORyROcJvIL5KV/1KmrhknRqFYEOHI0abgO2atGrrz34eJ+7M80iv+rMliieGBz1b2vkQtBP8vik
t2zlCzkbpajaYX+KMPjmBVa2kQBllyemkpvCK2TkXL7gqgx5RqGeFvTG4Jsq6opvax0HzQGFXmDM
04cE6/3/psi4nTa7fkLLl5ShKqIs46nSoNwBMLx2Ktv6xMkuZYdmT7nJ20meLwO1JocjnCnFSdVq
mUB4IWsI6Ehcd5lq985vW7KvOSGAqm89rwXlsCBZ8k8GBATzpaZ+IHF7anUWi+GmifRojrwg2Cb+
yAosVH3Jywoiwy2XzhUlfV8pb1bl+ZtqC97/vbvv0QUuJ9CnagXcC8kZLT+UgBWbeXon9HJg55Kf
iL1CnOcT4J5MAINOIhYJ0Xm5RbVfNcSypNAsKaAm2ZPdVQKpNjUWgVCxYJE+6nPDIY98FKWyI350
R+vUtc6cfj3q6TD1EPFlBEJq8fsBU9bdUBFWDEJKwYrCu1FKc07uktH2N8wSHXJSIpUvrbwAi+eZ
Y4j3VJxpFdqI5x75OcDhKeXG/VRR740DGR++tvX7cpLqWIn51g0JD0NNsoRZ1AY39/t+yxcK36j2
mPUUsPnI29UGlWOUMUcVWBCLUffrOrHRltGwuQUJk/2z3mtWmR3qKwK1Qfk1D8ShIe7KlSkgnuRe
f+i9pUXN42UcH660kqnONdUXsTT++PFzmD1EzCGRDkoYTmQkONCgwEz2PO3kn/F+eqJmZES5JGu3
D8KAqiVkrgYAa2hYZsEt5VJ7M9Hh1EoydiFS/j9/jBjg9HUdKWokGynRSbcXNcjiyC/1puk0Oyjw
HeCvYNTZTqPn31fJLVCoweQiZp9uLcpl6aBNxDkooJ4o9MsFDjquaCbgjkppwanfmYfAlEkwB8Ei
FsMbImm5KHi2dh1VjCbEtOqyp2T94eqzP/wlL0I3EFy2Tbi9/6Gkv0xCIrGP/HvI3xlwJNUGTwWO
9WUMtPndAAqBN4sDUHESgvbOAg4dUU73vquFLSJUo55RNpitNOTSXD31/0iplRuMnVO/bABDqm7+
c2TeDGz9EtExx3kuT3bVm5kmIvgye8dmmWBcNapmBlcnAVgosV0N0/hLJxQvMP81K+So9/AFZC59
HK9OWVXKLxiYUxDTtty3E7A549TTTjj4qSDcaWGxNiPfuuyhBHd7Ddsx2jX5pGUbNO9ZDZJJS9+c
qGCiIrLbx8YIOPv9p9VURWQ3uULuJI1xvph9ZzmzViNhNtB1x+ZnxCY2m61Hiowz7UKyDvOUO2lb
Pv7Jm/4lb1k5goixJtj9mmAhv2Ymr7w8gbik4iRT/EP9dQw3NNxOikMZKR9lhhFqQEWBRnw18R0q
LFATHs5zhN8Nq/+UBDX5TaH/ntKEXQBOgL83ZzUNx6+dPZlmHv2KRF2C6DsksVPeKgRssRMouYKK
F0hZxJ59CUlaloG51ge3zzGjrouC6yDtqGpgJ/3hWbYZI0nk8gu5fALhDmIqKLs4BPBagb1gtzNK
rG5hSxM8LJ0pVYBNj8/1iDvtv0xjsJrtzntdqEo3Av2uBmKnqdinGkSS0qEj6ULgDYkRjF7oHJ8L
aI2sJj9ZesrDtpHgWVAg4PZAP42BXJ/la1JbMnrSgPpHgxJk1s70QeL4pF+dZ9fCt8Kwzg/5joDE
I3ocirJ/m49K85urU+R1GOjDhHre7bXhLSt0qCrjsJ0eJ2adthjrycE8ep2papm5uSL5M2y7QAI9
5/FHLOJriPuqBrayj29yH9kqmq0SfE2U0XGdv3rPigU5DbBgMFjltAdvQiHa599uZ84sJFRI1EG3
vac1o3yalyf8ps61zLDWu62NUVcFrZCfyEX2ZNc6XbweV/Lot3eT6bH+YSQPuq2E0wMlG5HONwbZ
03dUHVG+VSLGuq1jxJEXz8aCji/BL9EUYsFfJX3dUznTLJESGqXwGxWbbuenLSaLiaLKoC1+aen4
RmyNDDt62ZnpatJDu9xYB8ByGcN9c1RDlyuVnP1y9c4NUMGcUn8Oocnho3gVLld2UPO4yeW/mnly
pKsxcr7CNX20rqnglzXvFV1erHuMzTvaSLZ/648hj5B7rtntK662GguW10EdSkF1OAlB+EXTJ6bp
f0OEXUI/DcXBr8YVLkmKUSpxdWZkQKYt/6ivxg47eRxKl7uJnBXHNc4tQNxQ1OBacEolfduTsadR
TQzIp/TxDB0at4dTMPDlHZtEDBkrgjVhef0Mu2vT5XUYCo8g/2FMpbyKKW7NGLLcfyj/MgWtnwCU
oZ+BaABeEh1JjhNlddNsFNknaxA4zE9FSX7Hcy1zW1Z/XUi1oDybiCLZ2Bjq/76OtjtyLDHZ9LmJ
idsxzCdPhNCPsGhhHVOZA9cxpDsvA3NPAgg+yMvuQozCD2oNv8WU9KS1j5pXfgD0Perr3zOIT3a5
rZiaXm5sx7Sy1pN2P8i2syxYFcN379TIQL61pnb2onMX6vOmV+nfFNDywVjQBHN+m2m+YbMY7spU
gaXca+YwCqjlsugQ206n16MhwW2yQ/L3k+NcOJIYt0mAnUiMQYOHtgav7GyhlbGZF9gG4hOTfMN7
muho6EEwEq+aSjztgwHnwc6qzQL4QkizIwZrhxKTN1qX8SbNLr3wMCoeMtwQgsUJwhR3w5VeLqZu
RWYUcvyODXK6/xMMx8l+/8u1b7f1fJnt2JBCmX3KEUpf/3isjGZrKKoyZfPKg1ltRXS2ZYHiHTUP
77zEs03lN2JAk1lZUdnZ1hlHHzK5ZAFiOv4Hg7HSrY0rMNnjKBB46lzGLoP6+pPwGLlV01V9nzOF
DtFMxtJsTYlR+s31vzy5/q+redj1IkcWQZRNGjDIPOg6413hQJ4/Q352cVTwGsd5YjXLKNs+Kqku
Oj5kLBe7cIjxFPtVEDcrHYJzzsQdppdIaunmFLChJq3k072p9dmHVG9FxaFXoSy0/x5uza5ReCAZ
Y7OYXbHXwDLvQU/ZO+y5crmJ1UYO425d66OjjsNYbhlklISi0P+ogj/v+Pzm6P0L7TRTcpFWXYSi
XPnCoc/Wk2NSPtIZgIstNTWGLv5Eh+sjKFU99b/9wD+jFG7dbmnNd4T1MnsCYEzje29F4sDp+m4O
VWkwCNGLeVJ5DhOiHOkUBIVH7rktusZtI+bs1sHLDFoHiDM75aw0s42YwhPjWqchU/xspQMbVTXt
ICLA8UODR57q8wPsHXHIeVzbhPzhxGqHkrdK4SqiojMWz+3zgiopIlPtijivm27p/1NRGrxQwrwv
2ox9je0A7pbHpSNicmCxoSx1z0gitlTFufuo0K6gbvAAWHxBC6l8PEZWwrhHaW/i6TXBgv0cd3lk
x2uU9w+jxzVRhnunN/J1eti+hoTVrOQcUqaceLBt4rb/LLvMcC591NApM2f0Nw+vZmNRb0bFFt6X
FhiFQ2nYEl1d6NxoIc/fn8slsm+dd0ESsH84RbVLm3TTyOEEg7UjM+Y6NhRxpK44SL8GpjjkkmKl
3ta5RtoZ95shUquaUMK9AgdldU+/xy957BQ0MhG2gY51+4/pF7g1ODet4N2hwMa0+DS9yoU0LgvN
u09q6s+pMJzQ5FVLbP91GnmIY6I6+00mtFEyC/UPtfzJtnVMgcpNUs4qaN2NAk2Nophctki4BBVC
QXW6FWMB/Xkhn36VQJcRIbV9ALDw2wzkQtwhextfXybEgS7Azzxi2OI9l+Lw98rYo/6VJKwmakcq
tbXklnEXciSYkCbhuS8IuMbpFVFNOrBqFMsTfeuVVdfsIfQQ+pQFhvUHME52FVK5uOYTHQAMphTf
k6lBPIFdO53vXmgHyTiwRJkz7W3FdZullE03/r22P6p8CsnFU7sC4ET8dCdmjfptN+xiREwrJmxR
wcXpdIcMBFOIiy0NrgJWXbbU8DvlQsTmcpTNt/lw0HFW8estMcqH5U8zzDFevara/+BNpsaUZqWi
SCmwdblcHzm24RBMPRAv1iAy8XKAZP3BHnu6m8ReUVLV/mRbhfFdbVAyAeHFr+ex7UzDOrbbm6k3
iZQvdS/NzPT2Mu9SKkY9RqXz72f+i2YtSauU6xd5Qx5fGrZPlKzOCHVmqi3+75WMqer5lrsTlYAN
Gv9bQxMvZOvkx4m2nwzdfcFRP9Qnb3zJWNM29tmIzWtga4dCnjR+m5CmVBCEnkQUXpfYuTJhMnLO
sN/Dg97DfNMFds2wPfoZO3rwp+q4/RwfRHSQFTUnrkIGluu5JF2fdy2ohxjjpBDAvxCyLxYvcYUo
YRMcxTne3iBv5DQuDNItYBQj1qjJTqzzVPgu1Jp0OfEYbuAa5+Nfu/jqEStSKl7HjdGH4ATyAbUc
3hOtiR0NspQsqHMp6ewU70D3BNaMHYf5ejtDBgXFXiVLZqDiL6CIYPO9TaeInVFLMoVIhZ1u3npL
iZ2tnRqNn1hrtputaa7IT6UNzNK1+CzgEvNFG1WaSuVsZKo1q5Fw8Enotjr/l024H/cRz22G0AZG
IU1uVzYtEwyF8aJM8+gQY/V3dig5RenWbVmkFm+S2KUNd5BYgOQzuJY0whseNTEyxNWcq+jZ/zUm
yEKBzC7yCKoZ+9FduLsxlrDBA8URZ3u75HUV6Ylvu0ceiDJ/shhsIA7bUgOZuEHAJbFjkjKv/yWs
W/cc5f34QnaPsImAbj3LEOFRdgL1WaQgb7TPlZEMyETuwTsV4Q49cx4l3dAzFX5fytFjE/zub0B1
8eZg2dGr1/h0N6q8HKFN+QvRCuBCKXQ2hOdmnpTcEPd+tJhcK8R6J/WduleGqNE88Oa9jKn5W6dE
y4OJ9fw+UsIgaq+hJgWqQekR9DBzFsJQlRy4xJqH3lQt2C+6jJssZ8erlDEXT1YLgNQ7BkM2QrcA
yRxdLU0y91+2qT3sFBOhbtk2xjKPB7hu9waUnmSKzbq48z7me8HwKL9mZqRi8XLEiHBOjUjAc1Ky
kl2NLkq/lhoh0xE6zKFEigAVbaCdvMx5ec06w2hNNLEE/a3/LJB13xNYPYzPdikCT1+fwyCxaf/2
QsraFFt38Ug2cFpGB4FxocsVh0u7bkf3RId3UxPYLJ+c6lNfXwCq4wjAIO2P0EC9p3Wld1gKjP+O
cwutLc4wwIpbnEmsG2aPAoQHqla1jeFxr/A53EchgXUW9d3SmaQdJJqnJCFtIWD7ZxiEQqQHF00C
IDAljfMv0AumjPnqNVbBdHZzccPfGHSFkYe9VSJ9S7CMt/78JUfvKzOpkWkVH+o1onw4WrfWgygR
nGT+QVS4iwIqmgGkbBk++lQNx3xhTXiXrADtYJ99vFJA12eQZg2z/ewNe17g8Pq7s4VRmth1UHEa
eO86FF0radEAB1MMeYk47DXUDbiBGIuw1WL2QQEP7vI5fDFo+Z5UCva239yfWo6C9k9EfaPnKKVj
N+yMtJqfTLCk8b6uC22mad9rEA9o83Qe2/DY7q7dnIsBf/VJVWOvx1XTbbYEUcf+CQnhQa9t/KoQ
8C9mlQ+U0wH/8zSBEa8C50/oss394PHo37EU/tUkkNycQai49oI3QGN1VqtyZvQ8aQanh2iQD06m
0hNCrS0QLo01gXuh9KMztSY6LR0iIh2m9Yo8vjxd0vrm4cT0dw4f+2rycA7Z+//pZyJeFIiJEdkB
MpYYI7oS6+snk0hfX79Hu8nF+iEnv72AEfiAtQmI1ZghL5D8uwyyACThYQDsCfFrwFDzzpUiQNZE
lp1Rz0HxK/1lNOnIeEdbF/YMw/3yVfzHMYvuN548R5m4RtqG4SDjmQaC1ZImWSCRB7aUI4yg5xMT
YBpZWJ8GavrsljufMcgx7+hA/4BUYWx7H5ldy4pTcmUqvYP2S38B2uNbQj7Sdo7hdytt2gXY7zQl
dOrUjAV5vYvYJzaOGhUZzbmIyNqvuvwsbzAQ7Bs2bxfWlR1uC+f3sjGUj/Zp46/mTLUj00aE+2bF
umAukvmHOurB/Sj93KNkfe0psPLT7Pu4iZORX9Z507g1ctciV1PpeB/BSqURxIZoK0jPemjHsaOZ
R3HEdDDpzKr1rZctWgbI5HFGK/fLKTbzw2hwOtno3/gSf/eL8oYw5eFkrPOGxKxuBNZWYern2DZu
Cq+eAB3spjTvz/ftPNKNuumpkt14SfwhurcAQdHM7Zo2c8Xt8/BKv+S1iavjZY8rWxAeV/mrWlc7
i/sGR9ShMtzFEtnO9QMayjAvnHgJRsn4/RqwkdwZT8u2JpTOqdf4z8UlVK1o/z581R8o6AyqFpUu
9lPl9mbb03obXHf7QP+VdqJr2NIx18NYxOqF7zNMMqiLP1e3mk8iMteeII8KJjGc/xWtstUiagry
fy6pGlj30PwBxXs4NFt7L3K9tZb0RmCeosJ/6Q8CkSTYbjy/YZLF7VxjY89xVWORMplLa4Y955vz
Jgkh2z6LzNPkLWz3YKGXzslrfD8qVaFYLh2ddaRN30T2j5ieba5V2rFDa3rJvR0QFuau15lqkB78
b6L3gfYa0aTqnnYxRrFxGcXkUfCmwbffIYxCo0kdjnRO5gmwP08jyes1f3q2dfpKosXKZsQohM1Q
IZ/J8FZpUJII/6lc9BXFrzZJMABi3QePm50I/UpnFRj2evRupDIYN2Gwprbd8c8VOrg2/t1VV63M
pG5ex51x+woDYk6DRg/Nr5OkZ6BRgQJPUMZBHXIQo4yGY3UDzgzFfC9tEA82qhRO5Hz7fsv8c96p
PxaipIi/t1VdyVCEOtbtJ0QKo+2uv15NMin50paHSwjjzRgevG08a4m5ddTcAFfz3geG/fYiTRm8
kFmpXxZZRCAdL/K4xCpFtxsRhASvau8eQOMgdMFWV2G7s9ad6L8nxqdi+2JS7Sb/TsqnXIPI8Vws
FkVBKGpJFD37OgAeXxF7tp40zNO2w14GPaLURjsWk44AXWWn9RXFHSHSVMAs4IZBcubJhc3cBO52
8x8GGkPqDkIKky0XhpJYxKWyUiu4G+qM8Ilme8lfFOkNkeY7kgkghi9Zu0eFEelOurVNgBN5g0p+
KREf1VABHlyBKrFPIXwlbL3cAQ8J3St9prGQNoi+CSA4DWlmhV8FDYypIE38J0mAoWx7rFwy+Mcy
S2/oLaHINuckQFlAs1w/JMzyWIlzYVwogpnWT6sMRFV4nQyzYCG5owRFAbHlDB4fNfgM+L8MIw+a
P9dRnMh6l+5IaOCguGtQoavCM52lfOaBYadoNWUniA+p8MGGGTmDPkJ3EhpJaf784JicwcKg47UA
cLnc5j33Ql+t7+xfMxUb1QJp358s+y/UJ4f8WhBr6Bgbfgo3mZFYC1iu8UShOmwmBGbITYQ609Kr
R9lLPXHoL5H1PR72AMSgW6v3rnysD1AwGYavTntWl1omCiR0YVMv6sHO1blV7y6/O/PQZonfY9jY
csI03T3a/WYILzEHEdw3CiOWIuw0mfqsqeh7yWVjPbgun0zpp1Tu4/U17MgidI2qF0PNzUIZYQkq
cnu8b0fulGcXFRSkbWPaitSdg0Pg5OoQx8CfRPXNEqCw9ceDJYB3Zb/MDBvzqAZx2C5JWFpZSolq
1SQwNY8wfBUmFRKZCBD1G9M+sdCb+WczvNg2Oo+gHSObT5wVsfWsNOvSmI0Zm3kWPk+QOaQ09Rmk
HvRitQbC2qgHaVetxNXX6bCJgEmfx4zaYtf3KA4eKywXvw6pImNwcckKXDmuWH9r5Nsk7a5S9Fmj
cBilXikm/RUBK9g4T5sg879ijf9NQYdmEzJm5/JkCLRJgGMJtJ30+SGewhMh0YGlvYWnrd4yLWE6
5n/wSVsRUSCKYfJR8yZj9YMc2puHKZjLgnTxGTniDiSOC0Tv8QKwaVvVjjmmMmY5qHX4J5B1TcHs
sjCaDp7KpJ8MOvAMRQ3bjsAsJbx4sfQUiQ1JENBtlwb63YNqh85kBXHkdz9rJnkWn+k6uwKINqKs
q4k29oPsmpBayDAji4iwJHkMKmsdSNEjM/SPayJ03htJdk27EkYc3jQQAE78XdyBDO5FT+zFvGVH
3c1d5hboAo4H8YpNQhzgd8QzkhJAo5v2+TEgNy3QikKht7rmgN5TQnilFcVDLTVgDfEeeP6GTCH5
rFb/r05Kzzg86tccn3yjbg9faM9GXc5NPu74irGvrsXM1Tjkb1xZ7AUgChsbcUf4Hcww8tb/uR4c
A4KH8PQJL7jKJF7ikpBvaqiyku0DyYk5ODrNnXPtjeG5Sa0mIIH4EERFlk58XqgIQEVC2Uf/9PFK
udRweTh8olII8fIEbDm7VMpn/BDyQJ1BatqUptYbQ8PgSQOeyujDx3E3Oag1wybh2ejQzN3XZ2Jh
Kv/PE93GvCqbw5Exns8MUjodbPFaXUhIgr4OhcmtJDqxW4qW6/Dltv7OcZXrLOrplw2gvDzMhoFU
scjWcHk+3McVOUWkLLG2taeL/wcsz/Z01CKY4SGtmak7IQnIaXjngOBeY5IMpiUBat7nilxXbns7
ryIUBd4Hqm0917M3rPMMY6EfK0WTDlA2czjATrwaCPzTxM0STh/UMtWqGvxflKjXP4BIt9nivWOE
pkET4SgW8AoO6S8IBITZVm6srftd0BXUuIzGWeOkEMH6LITubFOjJpFR7Pvt3hqiZuWjWCYqskWI
2k2IdhwMHGwlbIDiqPtfFJsgzhZ7UVpKW+GXGFBpXq6LJDzi0/jJS2kEPxp06CkHhtEXjbyEN19A
JaW6JGGokTMm37GM/ITQSDnNVAbjXQhxjsGZf0LtZiWsjKNqnnkMKuKYR9yi0B45FXelLlpwMZQw
qJ+ulbJdi9xERv/bbctMHnjow2OoqDiRBVXnkQPRUazKhONBvnS71DKP9F7Ph1x5YTGlqVvJdY0w
jbj4lqw2zU+QI32WloAHeKls/kkXhz1dmfBS3gYqCA1+lcGjF5bE/bqZmNuuzNnA79FSvGLZZiE6
29TjNhOBuSCE7RKqAbsGbJFNA+qpQc9oAB0O0gvS7n163SRYWGmjv+AO5LijowU3Z7/wLOgE7Obe
ShXy2qk62P9uCLeqhuclxPY874iVwRtx/HL3W3U1vnq7Hy8Fg5f2V7NDFaX6pn/BOMeAcCCkLpPV
kXGbtcU3EKv4WGQ94zK0JKbx7gDjfU44EpOc0I26McZwtezv4bvD5Vc5mGa2IjXbJDhw1hF94ipP
KSkd+eCPDAMtLDkuGH28IbC7C9nU0Z4y8OIDnooyxmx3z1fQdW0FKCMkoc9BovwG/t+v6AQyh6BM
j/Qr5CF8PjbWf2a8jLb9nb9KQRgZwXxYygqWmNMrABkxJdOc8V0Fo/1bowMAZNXxvgMsuFrCG/SE
4Ps81aeNvlQdL3ns4pvGVcbjBuBOU1YofMEUq1MbN0ELJPYYAiHgAVDnZO22qjOgw64kADAX7BAE
SS/mFghG4P/6nhQrmpltlZCrN0XZMCfQL5SxNz2YfsPkSBS6t4L4mQWG/pUA6Vdz0uULhBwy9jWJ
uQvrasfb19uaxu4VYTk9djNOZUuOEukw4CdljSSH419Lm5BD55NCTyoHRTKiIcEwQgEfD8sSA/nG
3wQreiH75vWdc8+EZ+PtHk9Hh+hRFJm3FSCHqv6xf5KiquO0gQ9+KG8jcxMCkasEwUp8P/dRrvAN
liW8NAi3ngvmrhPa2V4TSv9QcdTfio2QbFIUZLGnlf6LQPWTzZ33hZlZkgkWwOP89aSqhlfX4zx1
+4hY9M4osGlM6l1UzlivzorP+6zCb1FPiprT45JukrylLDwGGrWHDd0JmVxB7KLuI5LMV42xrCL1
KBvKEgMT1Jm47zw3Pl2QJMVASHDYO5Vxo8ZX+qnNJ+PuFe91q/KL4GssBN3dYQCu8zIyKEfwM+DD
8BFdvfryjuUaZbK8R2jrJ0RYol3cLRoFVpUX0OQ3XyKidRMMjyYcrDXIldgj8uUpFjORr0M2HUBs
eP49I7gpAdd0JenIPXSSdiNnFjPv2jAfDosbQVuAzHvWoLSVNC+8eqA6rySWrrHZO/xPnRxnwVW+
d8u/2F+oB8o0eAOHDcMddKSxiywXgwEbkoav4ieNnQepjFdYP7NxrTuAXAFo4DYKSWxuhqGEOCwy
wQWk9JLtnJSP+ksZKP9dVOrsGRZ4DAmkql64pCb0LKANyYZ3KWp+ojvZ0WCBXVhZNLcyvayQGpY+
jMicC3duxW/8iR55wde0EIfCDheTVaIfSHtEUrG8Z0mGZ24x+4G2VWnReTI7hNya5G2aIK1KujML
cpwISIxFvigbKsmYxCXYIntx3fgysAeercqsht/e2DqjRJU9NjB4o2uLnV5R1rXOBG7yPUpzgJsZ
h0C4Q23QaJLKAxxuOkQtYqHSTAzdz1z+tei1wFaGAwC0N9yViuOO870A1xGFtHnX7UvyWPcg9T6i
E6nHy20F1MkqYL6vNGlhhRe4dY2n+N3Ux/UmLEbxTLvRt1knaVAHO7o7HrLkHA2QH6S5xIG3S532
51H95gHxtDyl+Rm8PAkOimnqV7SpQmW/1mqoEIqUbYKj/Xg2rJ5PF4MaiK1WRnbOMaM2fgTcyTVp
NJYQlWaZ9kivLb8jdAiaVO+PVNpVLRFe9rWRw8bkrQMzaRo6S3oVJone9lT8XQLnwRJwyI217yrA
LC6WP/ia0kdg/YCP8lgCZ+i/GFQZiZgDZ5EJjAuUTpFfyaMIl2Z70reY9ZFtzynH9ii3AiBtLCLZ
njVBrgYcyqcyXwvBt6iQ2A9F+FI8FdOAIOSMNSc6jhDDfrP1myo5PGbKlSuoibkNbkVZWApgCaRK
QAxoj3mJl2zdmd9imInTEAdTQ/ZdOjb9YJYc/7bAW49UXq34szQOBFbZgzZymKesRQ152Y/KxFX7
kO6wiWVDa7sMpzu8tdL0sf9ktMFT6L4vg4c032UonbEnSgsjiUNxkjgWWR0FX7dkIOjB5mhVyUJp
Pu099Zg1cNZJNrz5y5adtmU59GtZAevayJmLrHp+j/Z0uaLPDjKZC3fPNeXd9TG+oFn/mIttKOiL
5nrsNgl1TRD6QgMOa6PO9Prkkw4aZP9uuAeDZyri3M4hmNma7qZ41M1Wiqc0NKdU18hygOvhP6fh
EVyUUprThHKN/VJnihrQ/edP2vah799T6SjvQC1DhheJeYFnr8GN5QV/bbcVjQ6C2IrUdoGvjjE0
ghDSZmvAljS9sS7c9aVhoLChaQgWJzlxvXl1FQX1coq35sRDsS3oWvneULlSkcIl7pKUds4Vo2iR
YaMyWZiTw6WxSyaLkSstlyxkBrhpCMDPihY/Sb+LsDgsxPPw0EuzH5R785qrb88i0uAnuNT5Y0w0
Ug7qNbnjAmCPVXDfphoZMbg9CRPgtftH9YLDQfYzcz0YU076IFVaxtuR6idTTwzPHZNhy1/OTOvJ
Ndz6a/nU7FB5E/cr/axIKLjKH0kLNqZ+DX1V0HL/y3UguGz0OV3PpbFRH4avEy5amfq9XrY9tZdP
ylWA//lCcxUEO8vXSWAjLLimSHmwuLfbU61cfEAtGJ+PRaulewLW9FESdVVRYCsh4i32VyxMzMaQ
gp/z6ryDleLg0d2Dcz4yKKvu7CCsGAkPPXLRp5X/ehBDvLwaZ+sXU4h+yAeepHdu0TQgK8TaQth4
D/Hjhbc8ddeE0zcvXod8hLbJ5DS96lqFxyWJnUjaKjrAZ9D2VHTFsgdRZQ7R641WugdCk+CcIXl9
6rZIkNFJRbcGeocMlKMCxWtZl32wkx2v1VBxfFNRPqVfZdbza8ai32iWOh5/Tt/mOdb88qUU3mJ+
g43JtceR9Fd9zPVraRpsAccl8STUGnxr0WKVfp1hee5HcPgDdKMUZTYhyye+TaWBzaCEHBnUWl2m
HgHh8Tlwvf5o69Z9q6GRWGqi6MXEdXcO/GK+VQ8+DH5ZVKALi2jLrSFkWXjvANg7oN+ijCkDtJd6
Jwj6kHnNNMCIXu28vzZRR47hvjjb9WrMpBwgCpV0mn5YPAYIQfWmtKVZWsp2qM761c3A9oMDwkwg
Pbil8JGnodSbMx8Yg0uca3DjOV7BD3+Nq62enhbubZn05TJ1RsA1ldOni7164izb3K00P2HLik3E
CXKiqseRCOb8vEnLl0Yh/V+eJ7CRGc0y64J4Z77VBndP+A2xb5cd/xrvQwQWVIjT0tV5Y/9pwRHU
KmZDlYIScxZ9lILjkLTbruxCh1WekHLd4xrU+i03pb2wQejW/6uWa+wnPna5zFreCi6wiirEEmpd
PlrYfuky10HLRuCghnYOp10zDm38CPHmjS3YjvkujKRHegWogrWqwgHmU5ELnUMkINRvP106Ct8E
RvLItuN0WiMINWHLV1FiloTkMBhodCsGcMr7lWBqgGafu6ze2VPNsY4ANH9GLF/QyVdugFdFaYym
JqVYNx00BmWYcLjABpTMuH4NUZ+hT9iyi6uBmJVHnrKVpqceAkmRe0GTAxsf6e1ptcJgnfat5HIN
+b86uYDTVpz3pcOqEFlWXTk2Ymlj07s7W5qiIJkQnjnCrY8J5HU6xLOUk0NWjDq522JkoREWFY0+
SqbnMxkRDja9CFKbdlQSypN3CYHI5MlH/IOlu0MmoMHNIbYlUYAzMipCZqCajcI9fkjDBzN3BU/y
HyauxhETL/1tyk5DJMF4Yj/ER01dGJqeUBCk5dTxEYmfqUF66X7uwnH/EqKEavFhPcc0mDOBcjUt
1AMXMC/YbWqv2t+3bbXf9BYO+MUuzZ/kTW44cVXtAH0dxAwe9BTR573bR7y6NOEHzxvaTJKXxuWH
FJIg9qHBmcmVw3zU8oenQgMpfRLnHHt8tARF2kw1z5dobWj+knHq6qE1e2j4ijHDJmNjsBZX/osl
LG6Tqagn+YI4a2qTgUiwZjQE1jR8Gg6Wn5RaI2dBcrPfGYCyIBLoqTEGaV4YjfLrI+CR1mFB2r52
WWElW1zUc4ZJT9sIjzw3IAIWFTafeCtjgwnzjLe2zIEl/KBSbYmmsu3QV5hIE0wto1iEKjzK9j0D
CFZWv5g+h3Yv5BAA3w7mDBT1R/c3r2kDRIBYrYD/PGSeFGzbFBNsCfK76LP9V5mkgtcw8Z/2SDIj
u7weZD5vL6hUna8D5XxPw/eEOAervR6qm1xtsmjo77sm5u0LQJU3hKFF3TRdFHo/L2hyfsmMlYWA
2GbUUTR9l5tOUY+6yalHt4e8Yuqx49LH/6tSL0OL9o1tz5KUgZrQlqZTjPh8cKXwVUr7iNMIbY0C
DBAe6ufhCfv8Y5crnC+9jUoHYI6PTh84lWGdzoOofea0v8A2CgF1fTeVNDoA8sgtNUfZYYX1NKwN
wK5lhBCn1IP42vBbDvJ8r6flg41kjop99GQGnxmMRdwbr2+scHlGXWtzzo34l3fiOTRkVUSqbrrX
RhrHtU+/ANYeLeM30WgrPxRo4BkqPPbPiWe/3Mif3lT3sT63zKRxIrgSlB5uDZBA3QJB1f9ibGIq
3tv5VK7qWXJmncUWEmVbxw/iAo6mO4u3MuXbnEqSWaTZ9gQbxD+6DBFbbunJeAIpLnb4kx+Fo4O8
tRIFEIk0ErkmZQTngN7XiMeZOTYD6drM8JEsRqLoXeY1Cy9dIiOwexrMOMmhO/eRw39/HFjGWcvP
WUF4uzb/7e3o4QWm3B6Trlrpc40bx1Z4v7JR0D3ban83ONpczaScUe71fA//ywZNECyysReFy1WB
x08ogCMTJN/WS9I8aiqsRg0yE+/azrbZczpntl+RmJM81jBOLPgO3AmV8/BB+eEO4ivciq9K9437
ZNX5lRJz0QwKkyOaeSK3LnQOA17uUwA+eChhycLPkJp3cnwJUw/GWhdZ2ELV9DZg2fV4iQjJp2/2
b3cCmBxj24O0GKdI1c9VKRXqLo66DbtgowQoystMtWQbNep/RER83EFKa7wN3DpQvZhNb0tKqnjI
pvvW57bP3r8XgDyqPW5XXMwnSV9aGOPUB21/RYE1QurXDjZAXaOsUY12j+rHN2tJpUD5zO3w5oMT
5xJ6D6/gyz8J0aNMQGUXeYZJFISlbQx40YdUxUy2fpHb2necDw5NKt4RwZZQJhCX08VAa0WkVsEn
o+Lx9AWMT6gibpS0DyBEf5DRKI7E0KeQhBrrnP6Sv1uz+xWoGLqUKPZVN0FfMUCO/c7s9KnK4SMt
ghrS78tYdD49InmFTfoF7ppr3bzsRGo5biJPsCDRTZdFN/WKxF4TsQbvDB3g3GGTa6Jag0fExNO6
cE5ikPQHi/vwGiSmJfQ35KjqMyNJEIDXvBAgRlyyCfeDj3LNV4tCz1qCcIyxl4I4vLmM6cjP1OW6
JWUbVaijOpu5mHkmhet+u0fQvsx+jEt63VIV4MRkCnjBWOMAPUABDx1pJ2pCGce9xEsoEBsGB7M9
ySTrvU1n5svz2/XVLQxR4qe3Ma8zoW3k7MrgxTD2WuebLQTygcEuFSxrjFbzE087jnH9qg1hI+FR
5lFeRldPZxmnbMSecOG3MdLAEkUWW31Oxprz728H9AZbekT9IguZra4olGFljpAOqsI17A/Ublqc
LY+sMROwPtxKmrTujmJsZW6oe80uTifzT7z65qHa31KW4JAyi92LxAEfM05CQ6racqkD+PMKZVcj
anX0cTAwGhTrDYjcK+Cem1HO1gvVFocvwk5qNP68yD1p3hp/ec0Q3wkWxOqRk5nY+JvTCHJ4OjaB
kAymgAzIahbSrWC1SwJrq+NzNpoPBSbIuSuhkJgHaxrkNHkufCB99MxqP4Dqje4VViiTBEh9fD5T
MbLV6NXOjIHs5U6+rdfLYD3sTQj0J5J2rxxwNbjrekJ0hwzMIDt/y4B6w44VR0IdsUWr4XmT5zE+
3rxZQ50CJvwOu4QMy+vnz25Y47nkgy29jWHCPlcgLAv494o/yzSXq5b61hpGjOIeQyeTkOHRjduD
74QaP4p5Hu80yAOOnAsmf603HeUwK9fFUyPQvrhukSV9zafspSNFrZH38fo7e8K5lpk89bzQZ1xu
rRpwCifUxG4cO0TxVOH328xZHo4NYAabsgFZmhNM2YOO141Ia1vnGFlZtwLmkX0j6YT1oVjoO8vq
PyOqevsG9zboLWheVGIK50QpnEO6sIE40eKe7q046SKgT5cPyrJtwH3ukYE0qVryx13rMXrTnBWz
PO6FhjnHnpQm7jXsXfsMukDqNKrx0oIRxyYVKE4m7k8FezZDaUTKySaLyHqT90zE+72AntDw68CE
OlCEsLOmDLJbfXXASP5i0iaIjUZzwRXMcFs5oBhjeKQiGukbeqgxyFL/4WMdPw/HsT0CjkJdxxA5
0mOhenz6NIy3Bv1ZaWaKkqxo4CseEVcNAFF1MA2w1W0TUypzG48J75zchGEZOTwMhbWvCN40jjlm
IS3ji+FibV1q2YET9HbyiXoMtYJYG2nsm9Ol+utAs1BVyfkScxTg3yMHgghtYz1b5pS1WHps8zQ8
ldghPamXx+Wv/LpOneq7bCnRV1Zw4v/6+mjcbCmG/HAEiad5QUSbzzwIiFeJTXHve5s2xPqRo0es
7BWie+iDh1f7/zqFhtxj+yWuukejBYN3hc0FUEAChMFzcJ4ZGp4lFa6aMHdQJ2yK1rbTGCPevuaS
RzlyIsIOZ4bF5Af96BDuGHBAzuSDt6S6IjpkB9cVouega5ETsaQ8xfrpz/i4hznbdcv7ImJ7jdU+
JGD2kOR/gQfYWp4o17qv5sO0yLTZJRoJ0hGASWsWtD+e+63RSJ+nwgD/ajOkOFzgs59C2SaRrb6Y
8h0Y3g2qfb/92WBUR3tQ2A3whx8u+kjrKKbGCEYjuB4Goa0wtaFAXcdducF+DCtPkz8Mc0isrPk7
fFnI5GOLgujrG0gvOnOaTeCYGlHqn9t+UUn0F/DxweCuVscDwlxp4s1gLHnox9BPN0YbIJJGUEbQ
Uu7lCOwkaok/CvMvX4uT17sJSxtKp6FuRwaQkFL0qmVyEJgjFxaj+SoqZB2C+hIkHyHL0N/5cDr6
crpIxZ0xMavW2gEOxLzeJYiX4vSNfabwFGKERXqtQLt4OjUoqY98oxlHLrE/fExwSWXngli7GYmh
mib0/C91bfkWDU2XVfUACj2DIDthVVRzugbBbMDlUijEFXhVOrWjw4J379z8VhSljTF+/+G3EL2G
oK/HsCbKRUET9p8GlJsqqPr2wg6odhrwhXaxZ/QEkLqjAqSyicbDcd3Nx6Cuin8s0/txu95BpSYV
pxB3yMs82Z1b9GsvID7VSNtFQ19N8r12Gr72VgRsRpkBB3bzoUg0aDJklNZcF7z+a1zp6BzJjf/A
Vhz1HcxCKx6BHTVSYEh+xOqKcp3f7SQYpgDRedsX6hZHnsaujJCTbuZ3S5wT3SdSJTtZRdeTkRGw
oUpSMZrGSxuCtMxz0Jj8GQ+2PyOYfiSJXxsv6r0r67TnnxeiZTkjUl3t1PZmGw4lQejDGYcYRg53
JXpUli60QmKwupMNzh6CDkXO5nMzeVjWuV5sEOZPaDYNT6+lDwXrAh4KePR6gZrsIgvrboS4M+KU
AUcWmSfE67hUMaZJpAYtmFRwlNgfGWhSXfXQBiMFWXZamXzavNwyDMplKVkdwf2dEIsyEVDtaVxH
K05Qe3S2Dqbsy+j7yFgZRMN+b4QiVT4CVcAyEvd0Tet1v0xt54dGItc2vZgI371gGu+ObpUo8oFB
b41od5l/aYRKOiO4dD9eoHJ7fIv7XTMtBIDP6li6A1nqxuVU6D+b+pjo8T9mbfP5O/BY59We51ZZ
lmUTx07HeVGUHqR2dm2DHOn+/pbwsb6zjTAD4SM+41Eb36TPr3UIINXh4KKHZmGOKJkHxrtFBLS2
xOSZnd0G4baJLx88CZ1dVvETTttaHh+KcedguxvoG9dzFRJ9gNLRVxMHHY1hFW0ZYgYtD9LNhDI0
wWJjC+P4VjvF4w+9qNtnI1+MOAYuw7Ys7kMzZ9BO9OYOMvzN8ehCsqoHUTnOFNZQJWbUvzV/+oKw
lT/fXZtYt68+GwN7g5Sbc8ywQhHetQI33X7rbQj7iNEDDvBpXfOG0YfkaeJvre9YKrR6QRxFcxUn
wSClhzLn69DD/mYnAKPS2ajtw7TBU5p8EJqohWBUMWt4rlcMkZp3iJdUyMK/Sicsmdpqh6wERsMy
ODB/sDgkInlg5FpUNpCHAVPlley9je/GA0IpKQHj1QffhwatpCjTnqjCKwSsdhYrRSGCcso65nHI
ZpuQGMBCe+Ohgl9j3rI52R6zKUp/T8zIYsfJVtF3UPQ1199ih0dmKU72u1+irFlAPlqXirQ3Impl
puT24rpu30k3n0ostQOU7zNa6ZC7qV7tOcPH8xZ1aIA0eRBNI7x9ZU/yD2h1s0yilGfGQOe71ShE
nMvJYSc2MHiAI6a+kz+BnMsTPJW4pm1cscLcS8IRzzGzWV1WYnDZkUer5uJWvf98GJkdna976p9V
Z27FLvIQYSt6PtD+w5/JHtvGE/y8XWKgsHHPAC1BN2+fKCcDZzkCk9j7DK/yBOfhRe2PcdnNYAl7
abhkA3wwB54ONkpmapeatJOIoRoUGQ2yJl/Fj68KxOqHSwaN4P37jI3ezqdmoanfIrevNr2u9d51
JgQoN+GqnAcPzX+Z6j1QqZEjA5Ma6AIhmpJSHPpCYXPENxkWTGisKdrD7io8gSwZTVpFXRw96rpn
OZ2fis6ZAanm7E+HqVfeuaJKLgTRQlM2cjlyyl8v6VyBGBUxlmGE9hl9DjNsajQERXZ731twhv/C
woCHdjPk4yrV7qEwWXHQTch8n8sr3xGO9y4M9mUFcuijvq5KAZStsBhK3HiMJ7Hc8BmHqHoLuMsP
Yh3pq2sypX7LYujk8ooJ3yW61518n/pCajMmpHB1PZx9FmXn9R5lijVSQb7K61YbTq1H3daoXThm
GO4vF2scYHkjJuVPYQn/bc/Jdg382LaoY+lMGbvWVudku7Wf4pBKZIGJ3S+cqkpi8MGbeYknnp5r
4q9sYbWEn6Dj+TfGar4MbJBPrFYQ6VjdQwtVK1+aOencTzzTkA//JWyyBZycUgDT4FWy9b1uIOn8
L6kpXArV3DrZ7QDA2Btt7E1K1xEHfR5w49xgO8omum3SVSN2WSXZpYji2Oh5jEB7wh8VvKQBJUOW
8MxY6atbXnCWR4NethGwW7hZLb1U3TBH/5kHhqpK1QI63CFPh6Wmc2aPOEdXwc635TEcDA2wBADe
sQ4dWATwT6OL8CVR5NfEA/9hNmbIQ4Oex3TZ9dDkxcFIoOJAB1vf3DHKeYBhMpxvF1uYe/hlWFAu
kDpuI2Lr6rIFHLqJU51QCwZGyyoHOrochFisTin74F0sfndcREQ7zgaBmqlPJIprXDhedgNFHxTI
fDBQzwXZdfAsbbrxJ/Oo/Q1X2puAdqePrgxLBFeF+UC0dGu4QVXiy7rpJXAvud0NvfN/OA2tXW1B
UjKJei9lle5FrjxRLH6HMArbjkF6BHS9zC+YfP0YPzv37KC+dBiemW1XGCLwaKgG4LNkYnIt2g0Z
W4ENdhxQqJRTzvGrpeEKM+KVJdQnxq/ozgOUS0XV6kF51qwkaYPTp03KqO8g0H7CdS0winQl4wXU
YEUvIwclMPC2eksYG516qkRKRjuvLdfIBya2NBEVtrgB+icogtnZAOFDpKzZBKupDj5Ot6qQm+3D
lmBecOQv1XIl8n1iFEebtaZ3o/MTeQD0PwNevqwluUDZv7OJGl8lUiWjoRjZc8LQF/R0McdS7oy0
c3VDyk0oSVcy0+/xSsruuQh+UFU9jhAcaCL8g/3APzRs/J/2xmvZODDlt5txiNY356EuULbBEz54
y0hdGJC7nXjvGzqNEwL94m5KRhgmUMWi1yvf1Df8FPcbgSv6ONOtD+/McFXl66xEbYJ4ZwVdpQa8
X4aC5n+8smjnsRSpyDn21GIlx/cWwKAXYr0YNpErU4qwc+opcNg6N3aEBxLZVnp5VtBEWZMEx6kK
b9kXO8B39FOEWcKbxxgzHwRpx3gfnP7KQs0Qa/pwsoI36JzxjfcZiMXZ2JYan7guAJ2rJ5RAah0o
x8MlU5uisI0pZU9y5K3lQVsQsgwyPLfQoBQDUVX41NleiCM5356QVY+932mmx9rLwnwntjGlaPHk
2kd5zlPUfSI6xwlnnfZsg+SKDyY50kjMZQiWWZ5pR3h00JNFZp18ExYxPVHEx3FatMLYfqOxf6oc
LCE6P9vFXvAfKYEDzwkVfX5FvLoNk1uK7vclyt23P+TkUmF2k0/okf+9zHHFYL5SE2jGW1VzvtKZ
Q7SmBYY3Ja6Uv3lgRpXnyMNaY1svXFV6bReuvvwN7iuxBZkXLxjhpnSrU1aoqCnxwXoGHMCjq9UT
rhqzboqzr/FOaOmf0OKQCexbW61TcK0NO7hfASsaHuEpFIwYygO5RCj9NbOWvyjfIno1G10eK/b7
LcYEBu8sE1w/L84tojBYDOaO00GFEctzkKnncCpt2Eq3QIoFgJut6clBAse6OnmYE01/52anYy0W
pACgcZvTyoordgoiYg2l2FHEAsV5xVnCH1We8MR7nIx3WttrObyO+MSIvBAb3J03aZLfa4sg3mmh
Xofd/CYcI0wmTSPKpzsELMmtQuF+b8VOfmjwloFwbn62RMwTrUDtGyTtQrxw4NNUpwiH4E6a0Pfx
vkR1MgKl77jme0ZKedOMdMREVsMqZSwRP9FLccmdOUR5wrCH0pTzQaBos89bK8zDLAItP9pU4Egl
4tbFzTq8sJ1mSHdnBgnWI2P43E873rYG/q8e2QS79rua5TlIqVOddiC+34qEt7k4oBUsl+05qz5t
OmdLr93dOEB3+rVIVztD3DId1FP+h8tfELM1R3OQJKOyIat5r3Drqn9q/Pf2x18UFMz82z6vcdPz
MuP44mC8RN7LsG0CEcSoIQbRUjuA+539gX4buxwlYqPX3CBXq4mqfVfvORNbAE5ZKJu+JeboNp2y
1N3kK7FzpycNRO+gm4E6eNB029/qVdOMnyuppgfCASX77eVZbnLNRTu+EZNJsnIxbk9/1AwRJ9he
VYKi/lTaCZL3A3+m00kCb2NvlPwlVfULlqWTef5T6o5Klp1t4/RHOE0OPHJ1FH9UZZn9/iEYzAXD
6P6fINYi/4j06v+q85gX9sv6iP4KQN83uFXvqmCPDbgrGJFx2Ev6Bq3RDNImuvqxdGkspWmUIqb0
4SWpbjM/1Ki9+yEGvISjOcPsCixhT74i0q4bcUBIqozT5tQMoRhydf8CEIP+Fd19ssgymZLlcSPc
QADPFtA73e/sIe9Fe3aylcfGfDWpV4JBh5oJCHwNAsGmeyofglPreKWa0Ifsalouw3IaWF77q9sM
63fxeXqRm3cxwSrdRWyXfQEU2y47TC8z0YIMWKRgGpEiIs5ZQ4s5FJkX4ZV4FebepP3mGrgYlGLe
x6PbdQSvhTMtALoKN8QnMY/yVTad/PkOWL27tp3UqLR+tmGwr8gsAzQfLOfQMxDu2oACuwYXGFKV
ZUH3PgBMgufL4VCuJyNdlBzjIzZWGCfrAZax+i8c5JxzY//XgJ/pVfbf5gfUDmDRVIsNE36lU/79
Tx+YTzo82/wkqX0aIjh0+4r7bvRl7a8fhg1tgspCSf6yoJnSmNXnBD+varoWVyeisr3JNl8Fi8pn
fz3bPYEmWtOFwi/4xAiL9LNjUvIOwWLkJTlpJUMBnXmQmTivdvL0j7re86XzwBRC8fDCQ96plMns
pMZrmriKhTHWcdRWWbnDoYf9HKiOekUq+A8sNKDeIoFmjgZJxl/Hcf66yBbpCLExxvZ3BOqOJxyh
A5tGOFJf62pC3Zv4RavHt5i8qw6ENKC9m4OVn81CcIFAQuyzHC4WeclOwLQKqcYya5JoZ08nU2qU
x039WskW2QBZjOgOYKZHjUxPGXUdevCCuKI7uTL/RBspf/VHGxG6qCfqzuDZyZORxKVlRh2h4U5i
9rkGTV/aRRUtIF91oXeyNOCeopKHVLahAp3UP0X0Onq/ne334JJPjOhZqb7FWw6+Dl0IN1v4ZFUA
soM8ZHRl8A7V2nQueXwUkQJVc2P6VVH4CdRw//g97kiDKt44eVoJ8Fod40DYs/1hGanKOVTKARHi
PBv6OiG6eaCsmNvyfDni/2+zy5JhpwCUyJAwSYlvtALFVmkYCFO5AvYiqTaaiZMPXBilQWt99hln
9HUVMEH/zrOtIAEpSwUfsl8P5rF2ji3W3oWGNf47Ho4BEs1Abu08aGZR8aaKBVUB2O1Hi9RC+RcQ
pYkgsj/wLz4v46TtI8a71OMqNA69v20oB9tAiDxpVWUSqtTSAIImXq5Aig4x61uSH8g/gMpZkhPh
FZVI9wPfrQrY4mkAAr+rlGv6Sqxkp1nP6fk1KKycqd6myVMihfr6g5PIMwiEPgiGIhSL68vStBLX
BDWAKEQe4NWtbnaZuerG2TwdJA94d3utdGrFt+up0N6Eld0Gb4SMZZ9G30pvXxlTwo9SvFyx/KNK
zOOKhEr9gwQQRI3cnNzEA0e9viV2dAKPGqcc2EDBZCAJ8LG1tUmnzN9leXizhSfXf/PN8Q8rYowa
GRizRM4WM9Rpndeu9e3XT69WaQKslDcc5RvVLTFgY5NF5WvOR61atZuoFN3cZzrA428Uxwg4fcQx
KTWOVDbx6Q0FEoJBBxYGgi8/nv5s+ISaNak8Dao+Kg8mJQJ/hKJdviCZ4VXT5m8n7wVTaNy8P8u3
5n+4eoN3TgrdB2Pi2CbjyVi8GkkmCSBWjxMi/0Fp1RVl3AfoGkmG/n+o3AGM+JmPJsco09ISZy9K
HYWySU7+/0H5Bm+BsL/o43W6V4LUipY/gwg2bbwNqkPx0dxYeSZqXzUvyiRM8l9MvFEQFyR18M5Y
FjmgCqjqera6SSk1cTyjI7Px4LLsdWJGMzWrjVhBOa2dXn8cYnT4+bcwpkUt+HOP5x+TcfIc40jh
i4G7kMkyQc3rJGYyQQdnlGokX7ijadjqXLjJEsDCufKwpliAvez/Fj5swTmIW7dX09Pz2Rqm0E0i
L56OZzVdpceLMgdfSvKbt1VgiRJ3t0A9SCLJKgTLghaFyKjxOqYG40tY+GGITjAOwIM4IMsocmaH
NTXiOKZqAee60g1Tyq6WD0rR/q3dUNXMoPQ7FAoKH4NhVojyuIsEFqNo+ROXCKdDGg0LGbDoLSWd
cxVCj3iDgdXGS8/gagbHEpP4tXlxZrN/4q+zgblHA4MY8o4PTRy602VKdFGzmIt5C+lZ4wPmN0aT
DzPX9+AslmH7Aa/PmdEIr78KSHOl6K7TKHfT/7LHEF1o6R0rof0bx8dXQuJjvyS0Dkss3+x8rLZU
T9/tDgvOsQd5vuguZZ/PuON0a+ABKKnJZFL0g53XND8V50lkr8+1/5/gJUeLBqazk4w+IkzjthPR
i3tmVEnRvDUgiWl2SE4RWyF2hDyrudCFxBayaiAUB3iS0ELMJXRtKiY8VmFC08RxpuFizTH+ovM+
c4U7yG6UPpJ+W+QHfehuPqXrO4Nv2St6CVDIvjs90KUlHFeVcFoE2NJrPj9XACfVAqnjos/BG+Tz
FU5qJzTwbrKxhVFwt3+9qvaAPOajR5rZqC3FAe+IVbhjEgCB9B2z2SgE05qw2A57IhnxIKTY8IX1
fy3nTIpd0BmCqdk0nsIyqX6XPPS8xAdoDYWgPN7hD85lgcrXXKidhLgqrnWNcz+EQ+egAjhnYVAJ
RjbBhIaDsidyvejc78QbwKVCZ8Y84jWBdhtamIQadAiLVNznGXTgE8axIV3hOuh+AsAxRaR6vPlL
ScOFqZQSysIa5G2iVCWkr7JWsT7z2l9Fq/X7YSzSYgEDjZIb336RbfaO3LEC6BhOGCDq5Himu0uN
9v7hFAtZ52Sa1zgdLy7hirkjqnig3v0DbYavQsNBFfWK9uWnkVuEJM+W59paBUcTQyKKGc2xDKfT
zht5bo54WcB9emMFbf5Cwl9H90ls+Z9dg4cn1nEqbOOOR5t0Zo6EUtSyf4BwQVmICk8JOneB4+2y
nj5FAgwdWQKzF4UQ30Wl9a7hy5Xz16P8VtN2BqjhUCSToRZuKKrgoHi6sk98okfL9zvqQR3fWTnQ
VWfqr7FcHvdN+lA8I/gOG2opfaptJfEUfxyODjLs4nB2eVnBQ1Qqsoq3B0LXljS1jmpnsWzQQjDX
6JK9Gn/fK8AvKGmvmkcOHW5ceKUAv/4+vppY8ntfpAr/DToGxbI7CqBxR5qroHXY0x9RzXEwzlwg
rUdMuMvkgABOq7nbQxwoiMNUCXAxsDKp8ZbqucmISEBZPYPKvjiseEoM/tG8gsRcxWFEZsfln/kQ
jPCvMi/wQq6oR65zt8SckF02XaM0xtM0OodWChe810Wxm5aRUlbJDK4s1ALtYxpYE7g9y1Qmcemb
euoEk6TbU1OJGwRQYZANuN/5rc7BPyydeNmsC6EQE7WB65YY9SZwzGmQg5bFcrNfISo+oVKql4M5
x7Tfi+3RPwsHjEHp/AGwVzOnkFp3Xu5Ugy1P/FMmOxNJ4uTSXR63vu6ZdCTby3owvDC1bbF3BDqO
YnyHy9zGVHg3Y7t7hgNltvvY1bpy7yIQNFumHczmLZ7QoIN/PTRyAJ2Lx8Uhqtt1uyoFaM6c6eJr
FrXlFurVt/JqU7wBuK5KTOn8FC3EsQF23MMcqC7D8cIOQE0vMWIagciXZ/bmrEkjG7CdKiwlIgrj
sN1HJJNfGA66vWY5IrkX8yfV0FFGPHdAAfoiItxSZMfVndZ9SEkMVUmUWGa6C1kj8UnaAsAWiOm8
cvb9jEb7qqeW7/h4sj/ax5s2WPHZak3enDPSNnigRJnIeAXFTV0enUsPMAjO0eeGH1eg0BYPCNmd
ddQD8TKirt7ma6kGXjSBxaRS+azHU//Bqr+rJvp2OstltE28JCR9d9kWYMDifgS9e7aAYwg9BwVf
+5fXIn33W/S92rjWP0/vd6tNmNS52wDq7cF/x8H1vZz3S9B5rG1eBRTZr86xRWiCZS7yG4uk6fAK
t1ibg62+nwO8iKZ7XSnA/ocOVy9hLZ1XPJyaQcFeXHpKmjV+DeGWv8sqJuWI5nM14HH3WRYDbmb+
WZzfE9tFOv+WuATy+bX/NwD9prcJynVzkLoXbsrDcsT5yf69wOenEqo6TtaAfjFVTjDYnDD2RuMN
jNyFvprCUt5nMmZX6KMsU9SyNlmmL1HaOI0KqJGmWngnEfYp+KNvOf+BG2EA+1SGVNHUCWAvq2dZ
9yG5x12Ij6JegFwkhM4BcqwSl8Xo9WVYwbzUdH8C1mkNA/ot0KsaombtTVC2/fH1i6yARU0rxjAG
HpMPrmc5iX+1Hk5k74aD95/JeYvW4dkHRKDacPciseei2Qc4rEuDvtbC62+wm/ZCn/pX/0DqZTWH
LZLE8xT1MESfbVmgfNio55orxjFU3woVLwrBiaIoNimjLgEKAU9yoC7YytffZbzUUfHUGcoxv54C
9srGhzxE37KNwjkXsZsy0rPsbq4Pu4sI8yqztgSyf1mHAUCkwxnur/CozEDCMEmlpDXDF1ADlYZB
Ekue9VM90GOSSZZNVh7ulzQ/Mfoa1SxkBpB2Ly9MXtlZjTNmgQJYr962bo13HmhY5npQqbL8nI8y
MPZ2YaHpf6cCoOkSIZosRopWIFqo4USR7uGiUoqZJg8c+Du0jjWjdjRIkLPGmjsffORJb3jddob9
GFYlK5kJ712qTknGWQ5g/oGCL/34o9s/HtJVV6xdtkIQ+UpOV7TUUt9v+V2dwmZNireeXng0f52P
WMznpY9qWe3angVLskupw7d+ecfIX/ULqRtK1ZGXe7qEGz5IuGP7t7w2jV7ChG4mjySdU6tf++iF
9SOJUmfj9PWQS3yOlZ5+jb+JrBs0Y9Kc5dFClC7M9a7iCbMW96pXdnOUV3tFxZgtIBFYX1f1Ny1m
hJOQtHWaT8uAjkRO/umMjAWkoOCiWWZdCMe40w740J0NqbphO77k4yKuE/autnkS5t3mUMU9fCgD
5u3sU1iZlkX4krq+rThA3gA2anFzFoUBIWPPlywd8wyhgZXW9aK3uUeWrBVd5y3hvafvcZBqLPQL
4GmvO6LnbR3y365NHzECb7bRpHf6dkMMzFbGIMhaOBTshFp64dzvJUR06MKk05N5utcK2KPxDlpO
0tTDbPWYXosPldRCA9/eRb87BlgplkOkurxBIUWaWjze+KbwxPKZ7EcZw2W2OnNsl56kcbMnhSxu
2iakyEgSAm1PImT6i7kCUoGGly6ZwhjOVRv5y763HyqZNg9eX0jWtxMQgL3LWv4WGX9QN1FFSLlJ
bQM0CipBXEqkhcUH5wtWab4ufNZKY0REwumc9H7heeOr3+03hezGGKl6eLPDYevXh4MCbZFzuNof
IDFQjPGcbxNVgYN2UP+uJsPxQHwBMHQK10+TG3rHrEl41YMnlgSCeVvNwcbC/dTOnR/BrdknXQky
Agj60q+br+p0dvUvZVgtyl5hTNrY8otGnoiKc6iRGhluMgF9ooLRJnFSKSSYxLhMc+30Uscef4FO
ueHtXOyixfcsbr3GYIgL6LAejEmoeU1fxONAmOOWCs7qB0Nqp3M6xTsBA4/VctLGWWAqnIQ130++
vQDCS/z0U9h0KTO2jAUrnOc1R7ef0MYqAkv/QEvDyKq88GG6L0WjutCT8YkrEJvis4lTqlJTm7qT
bX3Ca4xvUCIk8O2xyi3dstXvC9GjzB/9c7dBtM7OTiEsUg9Dy6smEcC6SaYhhKM4Ly75PKy6nlu2
R2wTybrfev/XTiMhl6ZUM5WEqPrgYhV0TAr5cfwEXRbVgqOw4wFXcROY7pLy7x/k+xNrsp+8XOTo
7AQIX8rasbJo0cyrlToKuXdzJS5tqhehSPnFWcpVhjwdHnk+hjRCzh97PxcM5STGWgyTnFPIsJU1
ZKq+fcdM2cziFso2tMowTyCMsqyVli4ymD4ED0Sa9uqXPTHFvdtF54Mkm2EG4l+YBkovIVF0MFlE
beNXrvOgTNIX8NEl6dzbzQrArkei7AilUaBwVf1ULTke62ir89ZLP1Z7SuICdSAhMZmMnNRl5F8D
ryr0j251aTUCRNC8aeNlrWk58Q5ZT0vAzYwdRMNT5Ax0M62wZSc5ZtgtzHwzmH5oLPEW9XN0GTal
uJLbxwjmVDXqRmMAovapcoc3BdngXXMsy43xWz31D1RUCFdRNHgMncK9AGH7JAztrT3/6Kwg2J/h
fPwBMeoPdO5hUYJtK6UBBXArFsFbMGEwh20sTTHiuYqC+VNmoFcBXMCI56W7HaTE5avKca6GUa3B
4MxkOgxaoXBZSZXpHl2O2CS+jKEcCqu8pEZBuOdcS9bwLn6Yj5Dltc6F6O1jGGM4KxidxZv0ch8a
GCWL0pQtnjTchGtyVYkPWTlTsZgteS/UW8bMuraJkpsZ7G2EP5nRPPzSols02oRFy2uBWY5YnAcb
mHS1L6ou/k9zg+D20Zgbpw8nCkZxtRuKnR/HF7s8v+M1tWGRap4W8ecwsooqi7Mj7j73P6QFizgb
q964gJ47lS+9RaUT+mn1eq2kNF4LWMQepihJnG7PZNafkhyWBHaWxhZJySh32/yUFvMyuVXsCbbb
kIBCXCT9A98czUqZ4xGZcR5Ampk2uT4z31qFdhcWYarHsKLCdoxuOLTDjN0wffPl5nLkUU5dtDqa
90VBA7VKCzbQzUGfyAm+ngVr4Ja2fMzITU7Dmb0YIvrXWwacqqPeOSaVu/TrezCgRNAwX5/yPaRX
wUp0o25pMViO/HysxUtsj0yRTJ0TQleKK/IQUK3/mhfBtEUTCEn2tQJ2O6oAmiNA5JMaA0ICeb7d
D1AAWOdlaChFOq0lQ63SnzqD+uVTr0yvGZ4KV0uIqCcJ8TWhsRq+cb65BpWbtMgqcFBEM7Bndo9w
5qfPuuOUVCV4mB1zpsCPshNDRm4uPGTesIhJxq5HZghOO2n/p4v8kI6Jm1f7hS38RAaI4InP9j+f
K1mAP4tHAYjehnFnsz6tvCw9witno2S93L8BYRamtS1gSP4ot1DuknrtVjX+iVH0iFRwTE3K16Xt
Yo4XtZ0vdceIbm5jhQzXk8oXtVQ15iQZ1zSV9i3TqcyQByfTFAW0ktQxffdnMwRHDgHn0UmOjqHf
TwdMNCcZ/RXpn+YprcmjJVJd0Ljvaqjbiu9szPz+1Q+jMNOFoX4s626M3WOz4CK0d1Gq2cKqJPF3
E6czA1I68llG9gekA7BaQldCevBfBjff06tNSZ5l2NrKnoCZJ0NEVLAzileEndJa0WTj4R1to4aW
gom9zkHXaRs3J+RkJIW1eGEGG+15uB6IsWcblN2xNo9Ek2SX0CKFOTbkvOV+9WaVbfXjIu5qYd/x
WrJeOqviqIt0CduJBfgQkJngIGvGmM7YmDxf98Hk4rCSoZ9qAKVQkVWxJ3ATP01sCoalRccNeHNt
7cZcfjkHe+VpUgkD4m5b0Dj2EqVuJB7IzM3OVDtKk+dyuNnw0ISWsj5/G5WwAZQZJ3YqRY01/bee
C7SRs5md1eBfoqp5F8JILaHTeKmye5f/+B3SQYXoMqL/OBVxMaK5KFauZAAV8zfK8fngGzMJbtiT
uXmmbBd10D8Lo/++pXQOVL5VxBjPMdhQg9C4EcVd9AEyoBG+qNjedI7uPJ0vHelw9gGRkkUOLbCp
EzbG0LADiozgqR942jtrEBfaZonzAf7W2SEzGK12lb+ge8FCkpbsA56mq89kMZsvNvjii26b18cB
0XWXG3HlRIqCXR38eIhvw9ghyfHaO2HjQFQJEhc8USMv708jdExaizIZOEQzQk2ZInt5aKg/hKdN
tMTjWqYZxhNXcs5wMu0Eby6F8EPhVko6gaIXW+eLf8Kv2AknL89x6KpfHotVpVkisliQGtfkwZ6O
5b/tm3LdRAscjBO6C8UKXVyFCUW7V7hbXn5HO0Lje0MHIf5O7L1mx8uoJylnguuA/t8PM+0WQ0TJ
PekT0/m/ODFqq2bZ69E4tgx4Bn1Ye/QSPOXLhlfKsDcHeZLCRYz2RX963eEYlWau/lHsiz6rtZ5b
TEtL/wr6MRUjl3gM6BwaMlZXB2L7z5FbxJVTi0xM1YSdMbHJQw+n3z21Lv8KMcTdtGwJUhHT48mB
JjGXNW8/yBh2burErJyG7poQzJonrz6dGV5v6QLtwqvLXkI4Tq0BZh5MZ5iOBcZV22tMB2jg4imF
34fr9cK6XxUuE1BKXzvUL+edwdmFUBB5mEdzJ9NwSSwcpvf3oaaafR6TbSfSZ/U/5bdAdbuS9Icn
3FXYs5wrSMP3OcQzdbc4PCtG/jRgzNj+srIlgE8Fsl8SE1Q0HMYZKYX2B8hGIlYlhXX+e22UjZxp
vdTB/355huNZfkEtMyLHecGf7977TtIi5sfhXbveIjG57p91A4nR6IiSKNaud4xG78JTlvgNsEk0
rSX9WfwckTuyLNGVclJ1FUjXdrhFj1oX5oKfWg4BhMtG3r1UtMnoVRrrml/l4W0hMNpOWt5aF+3H
gtsvY0ccass149pkY7DW/MLpbPd6+Q1O72Cp9AyTL5QK1JV74kZLG3Gz2QXhFwdoQbjoyElIhZpX
3DhAShcSLrG54V6FICC9wH5CWe37VSmHBdHVjcniAkWLD/3WUSZ/U+nA5aX3YxjTqubAfMVOjrBg
p1WZ8JTGLwFgBv5kSmYVgoxwPKRvDMNJD0rWej3bfs/33jjZcxrunX+rPPT0D/nmSE7ZV8gB2K+n
GdAM1hr7qevFPjZtgvJLi6Ta3ysHwysOV+P/94Lie7BeWLk5v/rz89hP7jAcP5eHT/3Of61N+VGe
W0/PjBexedsk1C5USnxeVEukDCHU/wUtedaM2OWVYhrhlQdAJZ3DjL/9/bJUqtH2zvePiXG1W+sz
46ZScbOB9ArXBbvUm6JdhY07AOqZIUJqNCpbGJksoRd64ZBWSP+GKDrcDAK7w9zq0PkJWFNraMXM
fq6QCWy/yOjyF5CDzb85AYmPK2xaBJ+la6cGuNulqG3WqqULxvVtnRBENCuBjGw6End/CR39kHg7
jeeuIlnZw0LZp8ferusC2B9+m9yWbpts5V1iMwBYMSe957VH2zffH2QhoAg+o1aLSznBIsYN5NGd
EroZG1xLgCwVzeGmzaPF8JdvP+nstQtl8++7EQO6wczQ/921KQi61M0hGscItwsSK/W1Cv2lEwat
9eweACc+wVUFQt7Aui0PD1y50MAi2DMAk762JvQmZyIEgPlGHeaej9ym8ZIwi6U4H2vVysQbCn+6
v5GWUZLIDIY1P4c0wKk+MJ9uoNOfVUPB5DInFnqywDdZRBCMndQPRzwgOUpPGTGJjeg2H+naITnI
X6aQS6aQrH3hr4JkQJVNxn2bs2wrHugXJPkibjvJLm2kewJ5UcoC2ijXvP6+6aqjL+Hb9tl6Drc9
+tHfiuOssW8pRX98SS68WMdlI5j0PGbKv22roL+97FOvGatIaTdKpKqGKYEyHDr9aq63ONpZ81pg
f+1YTmUxWQrBLCmOxXF+GPx6nPj7mW4MNW8l0D0VJmWYr26DD/cxrqEhvXGMaBZJUQfwkBafZTPJ
MPTEqD/1ofWQtBZorHysHkXUj08vP/198XfPETh4N5lHoKAD/G4s/ZBZSizY6hEPzuugbYdjqbdt
eBTv0BrSQOsYKoVLdy9oALOzalZH1X/jeyo2CBrgG0qwwRgRO6BnH9mfz94zCGlAceUUdHxdCcG2
6Wc2f+ycjvAG4RjSeYN1QLOYksZULSwuFfBFXQtb5PfYuJnr5QRro9L3haFwMcajg7NYiQm4loO1
AZKr+LYTO+nMAv1oKoPVucTOC4GNsS891uXm0q4ggb0vQzju7839iq6CSFnPdZ+DqWpvFVZCmdae
ABohVejmLPstxw+nzJKTJVeWHLS7FOAcMJtOdndW7sNyTwv8g/IdvLEgnoZJD+/3fdZB8yBU5Jbl
lMDAvwmWhdGIyHR8+Twweki7XtlunYvkm+n4IW6x/HhKU1j8iNdK1MiNVb9CRGg/u2VcPKGjks1O
BDZwMPmSp8ejiOHZfaY4fcMdvKUUGyKeBAw9HyI+K3VBpsUFj18OtTaLY405DMMi9WdCi6ChiEFB
SEiJ/HDjlR4vHAurdjPPTbJRsU06+ieYKFjLVJoHUhMx19T/yWDKmrJArUM0wCWGQKfIiULoeGQp
fayZneOR3L42kxeInW9eXtDcL7Uqf7HKMjQcGu3nNPgdtN0eoql7iZWH+qWeDPJ3G4uxIVXBzrJD
ffj5JJX3IxEIME5QUuOnHtrbyCMXY8b3vxbZfMdhK1T82N2X7Tyt0O7FqmlrSKpAQkUkkvgrQfZ5
hlbI3EpCNI9jut5/qYZRZgsGwUn3URKLJt/7DQyip5SlPmnFA+F0cr/jdyTpVu/BUlCv6/jbMD+7
tqNWaIeFrPAU9a3VI9U2THT8470sA10C5HoveXYE+A86Et9cbmLzbEQiffdc4GXi7dll9q9GdXtQ
NuGHez/cA0CeBxqTmh1JYkovFPEdzbCJ9gWHCnilHUnKBEXYs0NcChgnp5pCxnuh0SVpDHXH3stz
oEj4rjHlpluKmrWcVeT0JY6bu3KHPK6a+cJcbNoY4yjWXnHoPTPRV/nWxM/BKPYpKJAGoSNkVDEi
hyoZsXjo27dqUuvyxseZuNcb/ybnu5Qg9oc9gtcx2vjisqLUWwgvk1cIccqkasLuCytGFL8WZ/nw
vcsWcUrQZz90d6iyQjhSa/4s9U7KEQo2jhEaQB5Nb26kE6aP+1B+RZZGzH6MBUvkNBwdfwaI/yz7
R3u6u0LVzVoJt+2ZGRCEw/XjYM/BN4ND6lgV4iwmVEovplUYlMtToOQ4D9g5j4NKXxw45MT/oenj
T83uIBsEFr+fvvwYjBEUZdth2Tjt6onrTBsGgXmBf3lxFSpEYL4iJzAy9KtJeY4uC3sG33UCvExC
FePWnv2nSTZE6HqhYhWoTadJsr89M3ookDRU1cChWj9CPcOisIc0rUX8kSyh3oxR0oOh+9sVZHos
fmaDAI7YxJ5vFQxJ0Thkyyv+W9vAOoX4fp4I467mfKsIrVbJBvChUMrXvAvcaNmnLWtluLLjdZjU
biWDrZ4fglvk+BrS3B2U27OurylBkzgrzPoa+DdmYt20RJXVgjh3rtXzWjdJ4toXswHQP8DRVhnp
7OQxeC7MYd0jx9JABzbgaaXhF7EIn1WW+p/vddLv/3PKD46dL6L2NcLu2817Q1lvuuRJSMP1K83M
RYjJjTgGs23bz5M3tpp640JMFSG4W0GJkQCmOaFj5QAHzLDS3EzO+MiZNt+NtuDQb9CHzRRfyaU3
7D2IRLXjzaVtUkjPSLQXUWFQws/EE3ZLOhNTFWsToR8TB0cEmbqcdjgH72GAC6aBn8vHdUScK9oU
IqQMO9ECu57hFP4XQ6fnalJUuiahdFSfULt5Da4bko2BsASnxMo1YwvUeU3CSJ9z/AQjPLruYJGL
GS5ZSl+1vOnXGEQpzuvOlwRYm5djZF53U0bRTPnqgCk7SjvtsT1o4kYiiBao5PMufiUPiP8VisxX
0Ec9dZi5UpVoq6zRWdYx2Z+0Q7qn5vGbsXfFCTeeOjReZdN3xhFgKEbOdGyE87QdDSvcKSHBSiA+
AB7Tth9GeoZTTVGoStwvdUsk6WNA9DNG20ypNfQnfEhAcfvEVszIF3zYkOhudnlAa29JB3lYqNFx
Lshs3EfppBY/PM1SM+mJGHOhtSdyvqvj+iWTPHPJkGI0iuHx+mQKQg8WO/nOSDPSNIKc/nOXsisC
jJOCk52jbltzkARp+n7OQaB6MxbCGP9/iWDNEzAGGEXTFDzu1rBGoPR+Rj93yrBCEfx2CotqUlE+
gN76EbjYLuEpdeN1q1Je6OlgP4Imnq+L54u9JvnNK7wsFVBZWboCYEWg2DuU8prI8Xc7UsZlMjBF
Rt5z6qO/T0rv6NUnuuM0bpN+wpOVnQ7x4He+p1IqFOvAHfCjMMLjBSmwc9ovc406J3G0HrjKi8fM
DOpxmoO3N3W/VS5p8aZuUII+dO1EfgpiEG+C/wBRxhy+od8prlPy7Snznv2T0m0acqPziCzNiH8M
GH0iewgPt77EPqBsfK4NfocweLwN2rW/9hhhFVfuRLbQKO8RpCGQy4KDZEgdBhT7fBA66Z6TcDA8
VWzfqg3OvQZHc33i4bwE/SefUzn4WSOUrFkprwZqno+0iSJjtWyq0HDsgiVgaiB7khzIQeE46sOB
bTfAkzM1fToUoduDIsNfHKAwRS+ZO+B4fHP2Gvl189RB580m/fWWcfWq6O7uMSpv/O0PISYVTx/x
KwaJFxTRTIBHay4oyUtu300g3JEGIy2IwEuQgkQrQkhFvDhrpMYKgWVFiLlEqH0D0y4B1+900srZ
53ek8uvAIcPKfTq2d5CDafiHLsDzjrpcDoHRCK/DuKspWzdYr8sO4GLH7v7LBnmPXBPKcWgHOfqI
7htIDsIE0ipgqcRCD+20OIpQro0AlDjBdOJQ0tFHsrSMyvaU0njE43V0mCXlEKxBjbwG4yqDORgJ
3yL67gZpoM5PTkYD0AoQJikwRvExVIhdqdY7SaSsMtve2TimlZsXkytmlhX5OfPQlAli60jsEaES
CABhaKVg/nl/Ddlk50VQwY0/kJ2Xje09dGu9hPGewIdTAT6iPJCLOd8B6z4Ogi3w/LgLO9lmhJ2k
+rpdjpZnYPeNDblzqThyY0S2sgG/8DFZY+r6stb8eTZ4k9ITAfG/0mzUe94405XhBTqsrUoEd9ao
tlQh0oAaG03IwozamxYubDovHYrcWOWZ+zk2IigZTsEgBzmVRGRqPgqTBEfNF77+KKyGpUd4IyIh
rE695dJJUXvMwZEMyHRH+RW+TrqRMbsgAUfNwHlBwama3kUrDozskCT/mQLvdSdkgNR+u/71elIM
aTwnatqKCbQoQeW/BOZ3DlgcI5qBvcELfcjkZzoDksCMhxIjQ5v2Lt1hAsy1qz7MliJYbqR9yO2F
WYbL6VVelcnCzVUGsq6akd58Tdm8LO0+J/VCept53LkCcqc6+8JNHgruSNsBxZHQrJFVYa/BiWE2
u9lyTXOK7agH+IyCvO6tjuB9tZ+Or63hh8bQQg2pN4WS3U9dUQO2RxkUqg1NxThlOci1Qqx6aMUR
cFbD9yACXHgzt0CzRcCj58XD9cioD1Q1zVUnJZSHaKwEXQn19uLKfwgbPyS21GJu7mSs0p3Se7km
1BKJfKgMNEZZzRkshB/YIp9Iccs7sETmvBz4n9XGEc4EgBvNJZ13MvfHWX5LFmaBhfidWEpdt5Bt
62lTzbKmDyz/QeU25zxVYZnrJh/kG2+fnjForJMtaJS7LLojRRt2C+AsOscgi6oTwfzIVUHfdY1u
uzmZ10mLeXjQdGVRgOcog5coVoZ+rox2/hPl3r3yxm/xgcL5BpM9MaCmlI/chAUSXqi4iiW6z1yD
ZGp3EH0R/Xc2R+wvwNUpdyIXrNn5ESiKoRfNGXUZFlgGXsS9qxav2QJZsX/+cb9hFTi94GJ0H1Vd
TwumacI9GEO4bufKqeKfRgBe/DWbRblIbzqsAVVbIfNeFEV6MgYYT2JZJBOO9WKwuMZ2adecAX01
CvokLzZ+7zB5KdUEAMEX8nOp/1Qbm5v6lAYwgkS056NgDQuSfZwSNpNZ+etFp/ec7HTYZmfgYTd0
BJ+MNHEirgjkstpdZ2AVIc1T+dnotwQo673Y9w5XuJdfUjH/FF8BG2L0A0YPcRsZoLLq8YttKyh2
7l9kRuOochK7UwXIyVGeDyw246s6/39ofLh1RyiAkz3eLlMYDQ4TmtyVs+CNddhfj5N78CO3pI+c
kYHOgUGjdBwM9EbdsPQGLCRQ6tdtDpgx8LZbbm1scOwPvlptcj2IvGbUSts3vaIdWZ74KR8FPibf
CJkjgeizIZ9FVL7EBwL5W8Xcfp1Be9jLiqz5Z9GuZAJU0Aa0HXRQkD6YByuOKnEwINdrzFf1Ejoz
NrXKqpmb3MzWSkD7mjmHB5R8M8dImG6MMkI3eVAPtwTvMTutgtvFja5sRAirIWHqylnwVxmcQ74a
uPtjyBpR6Ok3oskkvMjnBF4Y6tjbvhNRJ19zTEvMW8mXB4lmlskmXzX22JOVyNItPgbWGlWvvu5o
F0XXCruJPiFUEfo8ZxzfCMhfBwUsQYJ+TXBq3RarJDL1TxgsJ8O4YxmjYPcDTFanXRD/0Cnf/AQH
ca5rydt09WX5o1+FnSHpG67KodcBhSmO1Ab6heoYzMzOupSiS6xFjuiRSaxJhpcogcBKsHNqwssr
eO60xD4e13vQSGTs9fykulQhXCjJ1ib9LzrUvBZ0fWwrr8gVoLQ94U4afodqHsGK0hFqoKxTqZIE
TUThysAdUyyHWXKGbvPHByJ5/R4DUNMuwHBUGrkkHABu6pZEfRpr8zIIdJz7CqlcrSiZWwK0ZApQ
gFhku8um6IzRNoiN5IWKw5WR8k9TOMhd7BrHbU6CILYYSkw50UomOXSShK4pvzUviRiSRk5xFgib
id7HdxWR/elLRsGu8GSvg/fekZgEP5x5anHQ7UFRUX/xXYu8dw2YUo3HLk18At9JPBVqKmTB3/R1
ZQTKUXnYbQrMNr6fF/O+Xi7vPVB1GBzgd/YWLzbmy9FB3q2srhRy7Ag6v34hLSQ905nhkfHZMuUA
coKTC2yi++yyrRTgAF2bvXlKtUHgqJ1qC12ufwjCq1G0gtEDexUT13h0azMO1H9eXXSJZxpyAZPK
3JdDeeHvR1yFr+J/qVJkPcCB5Tf3Gd6QynZ0mSlqL5GeSo1b0B+bT1m1b9QZOM3rYYI2yiP/o79g
+B72JjvZ2IkE83s8e84lBPVqevWZT3aR/AHc70qKwwbL+bnlk5GLtH2BB3pxmPNdApIunSmIkrBn
M7ADsuee28o0rGiuYslsIbU6kdd1ujN3UQwuqW626B5MyPMGLoStGCN9arOrsI7Nv5gmyt6jXiox
fXkrwdx2Yl8sJEhbrhSG73YaTS3bOi1Nds5btXSul4qpURtsGFK1mwTt46jCMUxJxqAXP/isPgOc
Hgt/fUuvsJ8TMNUeapQ0YGF/80bjJhX67xyjNvK5f/xPGi7cbBt+acpyRxOL4yv2/uuT28DARHmB
TCRvISyF7Hv9m3v4O63k92t9PHx/GpNO2eI05LlD/XoT+FphhyEeZa8hVWtT3ojE3x06TdtiT2NX
FjCXYs+ZHxffOVRVY+4XkVWHI/+DukJVIaCFULrbJES/TziljZp3KjRsXoINcYG8f2VURhNn05DQ
uO2UPcDtJmJD05dCIh8dZ2wgjOGErOMUkCvZ3Y64p4opY2KFJUGRI27IZ2aLRLdmqO5HP/kQzTuS
82AiIHRzyoqQ9xXSjMaZu7YhcgIRwmNqBz2vy9AVDrCVzt4jWis3WbhcFB5mjW2hsDIRJA1DDWsJ
af+HVCFTIWdQ+C62iqHuH4GgeSb7hZTbM+fKAGREQJ+i+5JMxwiJvSdf2OXJAewP/BydPsLSf9Bl
6KBcnEQVv6v8AeFmMr0XOiPY4iJn5NImNm4RMsHu5HaF/gYInPfNyB8WFt6m4gU2R9kpUKDjN+eN
jki49k/oLusbicepbhN6ygJ0Mv+Yipgts8vAcdEiIJM5WufcNbGUs2kxlbl+IcQc68zYYdTn5YQj
ULhdV5ACA0QjZA8kjVk5K2DW6CYvABybxVtIzzjQHbYEFWhoZkaZeWChnj6gopIK9k8BSA4jaIXg
3+v+b2h8yPLn1VWUR8a/SdipR5tbckNrG3OS1cVLsqd2EfmbeN+JljQkY4WFSo1ukruGsn2nCedR
K+DqDLiVCS6KfKRscSgjs3Aotdy1liM7Y59ohvjZAM+ErET9UD8c/IOcwMgiQ09aWCTFlcxJuQAP
IytiMDevGLHSdDBFAF9abhRRgTUKy9OlhtgQzwaEyGhZTGQwCIgDw+P4U92M9vXYNj+NLJPoJirS
8S7gZSSVaM5QEEqr2kjjQnpl641sRe78N0v54KwPj5uINST/PzwW+vMU4XAGI+YDpeGofavm2GW1
4qBWF9MxGv4rCMB5gFHQWT+z3seoCF3oiDXgZm7ADOWOz89+7IxuFWWGqx/YS30dQmgAck3o/ms1
T0lbqWyOYSIY/GlWrx06Alt8PPJZE2QTurlm2rfU/J2hTvLxL6oSHaUTk2Byft7qMLRwI8t9+Ke3
C1t48UYarnqekn5xJAV0JMZYah4mOL39a1NRGhDbS9ukJWoeeVsHXnv0mL0d/KX8dpa/cNIVpRKT
EPrWMPfhPyD9kLeXPyAr03le3yFsHuCHDwsYcXkVNLHxsboobTiPYOcDISW0CaxPggwLaZ9Anl0H
uOOfYDXiz9AqBCyYvKQMJ5PKC62jSUSxOqUoKGmFfBgcaMR5hXSbzKh0Whz5Zns+TW5gvvua9AWl
ecHNy0xQW6qW5vpiBi/iWi5SBbzk5FrUKYtUsf8RhUvnsCvXMDRznHyqjycDIPFBauBZNec8b4Ui
zJomE1ijDxrxSHBFUbiU0C6XuATHK6tQiUw4ZJM2ZN2HwXMyy/oXBiviVel1k7/BBNshzZxmLRXK
aW0P6Iq6hsmCOLX6ZvZvbHbwid7VlxjeZLsnTLYPWcd7oHQbjdwmeEbakqZKjYOkYBb2HS5bgEvY
mXJSzNYsYbhbMf6TxbwaSanGzxGuYsKX/V/GTTgEhMVRK0JoPb0h/C/re+FMardeDmKdwFtnqIEQ
ZBYICuh9IGbs3xjCkDpdfyczZHeY9DEMUx0DuyzWvYFyuPal+c/p0AOEpXtroMfkcZSAjroT0OwU
riWMuBDLkAINp1m8lGx/Tssn+IYyBNaxgrXC8Jr26pHXcwhiTPRzRrf81iVbzG48Qcw+2AqNCxU3
oRY1TRfBCVHbFhCOF91y6qkeYIXKjaNc1sBqZ/H/nOYl9GP7lE594pMgWZCvsJP+lA/rVR8FZ3YB
Q5gButuh/jYlW+9ZBQ+j7epZzmu0gLFwKbTa4yrSFRvo6YN2g4/AWxeTQFAZDq024T/JwRXNZSZI
7mqb/aO0p2haSddm7ev8mk4ucWODmRgX9svBroGNtMJhQegacIPaxL0dA7xriR3Ciw3FtOEzI3Tj
hfnCusuGqOgAJFPGcDrTANY6I9CnhkXZ+Ar7HeviFuJdr+aeH5si8FlxMPpiKZLH3wbAHBO88Tyo
a30StByG+vjeWsFWBmzHw68K0icFDfwa+Me4xZjUp+l79KrV4cYDTrSmcAs6LSu+jvwVKcGUMsQb
nv+pIsNv/lDohmO6DuyClVmdARQlT2rpu5MVmFtmsKYJFUfeA2m6L1PziWErq7Iy0EQ93Fv53U7J
txkJF4HToRIodLzPnwbZ9zUGsPCC2wYcdKXv+u013TLF1nRH/Es4oSMsKEpiLlXbi810dnyYklqT
e5nTYKb7g9S3qMDHibti8MkZdV+OmOLwLQs3CzDwoDu6/FaTU3n3EoDxvV0ebWDL+3OSEkwpUjqO
k+6YzHbuHqleD7fCf8hRZ/+mgXV70kF3NDxBJfKY2s5A0FQpTzNIXrbAkvdjyJ1NJSFa7WPldTrg
meNOoQr1s3hu6OFL4PkKHYHMY8r+HSl+I2BPWpNdIGVJ07h6VOvNL6/gNwbC9scA0nYlTlLQX4+s
CLjxtKS2s7bOVeqQdFr6oEvz+oqCVSLz49MFh4Yss2Z97f2R4DU2xpDm/7PkbuJWnafo8g3NKWSF
Mq4Pua0xklpW+VdG7qV0IK685G7fUe9nfPTYSjD8W87hK7O7F4lFNmtd+8UpKERlLzOQvn/a96a+
7xDd4qe0jtvjuB87VzqbDTUlyhHoAT/aD/DvRP1LrXqWm/ja1lbuzHf5DrRvkJPUABUdFQ4NYDC3
j6zLNRPdC8LHf2bNF29pz/sl8NgBA5g1xB1O+x217B4y/vKY6xHACMhELUcYyCPMAhf4mOkXI/CL
rDbCe7h0rlago6ZG/IMgp2BmQ8QwjXQ5V7/HmQET4kO49xysPId3JoGmZKV06UbPFWMlLirDhpvI
ojmDVtOlpBrSOxR0OwWj5IQc2V4iYK4K454zu+X8mskLnEcIjkFBK8R0QOBD7weLeY4zCqULXZU7
uVA7aF78SuIuSyhqnEFRDvYcgaxMe2QYAeGR5rbNuxGCz5wbapEtIfbQ0VMX1VQmGSaxAzr9vu3S
9sMG8be2qTUJialAej8C1Q/h3cGvdIYJbZGYbHp9XGriutmmZE9Y6iqPn5ivUYRisTFJuL6g5uWK
hwkxRW1BwTLVXiZZvthwBZqMNIWClGiX9fwjsS0xsNslyMaXVos4UgWK1PYxwHbGn+846mJrkwRH
19tymu9yLo/ANa9guDZmQuNJlezaQP2UXXGPYE7ixA54ekrdZOOVV1bpBJYHjTVDvBjyt3AcSPqL
79Ou+EDsmfmnzOzjJRU9IIKnOjstWWxDBhnAoQuYsLFHVhsMefT15jQTdb7GYuqEO7uCzIGMm0j9
JW+yPy4Uhtvxnl4g8R/2OAfeM0ME2K3AOEYQnNAwYwYfcThEZMHjAcAqpVWVCgSRqMufyMdgjhOw
vDpDDzJYfwfXyxvPiSSA3qB2GyXl3TLz9RIC5IBiinKeSDAVoht8Wh360DbIXxcpu+OsLLHDpF9m
41eH0NjFpGRrm1dxoSq7nXaMVCIu8mPPQeaiQPdHw3kbrcxQ7b33XS4JwNBAF8ONR+0IRa+Bo2hB
yWTQwFRixqvBMAKzPgfkw3IEWF0o7IjnOIUyiJiHaIjirzrj+g3zcgGtFt758cpHb8DVR8i+OV0i
w35jZtBGRxPs478KzC3Dl0LA4dnbRP23Jjgroxicrh3Ek0VOlBMINkuqEak0KmKoWT2oc9TRAaTv
H2nikO9Tp+dTNTaJWNzjB2YGVM3mjJdvjM72LLBw4taLMdHk5AsALvDOXr8ddcY7yYUH1DUy8vt5
6lLlDZES7LEGEorQ4sPE6JarNcpG7vhRby+ue2wJZHFjKF9St9E+QmvgA15GMnvmOva1hN875I4X
PZxKeC8vRWyE1MMPNZf8rIjYnM18ZWdO0234sV/QQZDS3v/WpKcKG+00x92zwu5MSAopVO/amkUR
fylXqT+bZ12Y4Q+OxdEoQkTMtEzymsABFhe0m1uWlGRHBMNcHK9CTeKNPr/4VTMkKrW2uUBCvETJ
MTnNnzO4N9gwrBA8LI0fnFxltyFH/jjauRXqRt00oaVLkdROoXn0h+FlY5Xi0lpCV7M1mEZhJyUo
9YpL96GDayT9CJbpg5hWg73XBTs0bSQJfFHv8PvfTmmO4qsG3SnVz/E+7+oHzeKZep3pPQe0Djkt
mdUCGE+K7JSeUXEcsG2QygLLyUjCdzndrksahoT+fiiKEEVw6RKS4c7/TfRB7jAH9FcE5ikVVCjR
3coSBO0PS856Ko9EkfZXjIZuZG2RO0I1mQCU3Nxdo5hDvnuMWrSmxne5yXOGLsIvgTGY/Z3wItqS
fY8EtDEa3QC8sJXu+tO04JLpaF45rvkP3K8d8k9WH0RomgTwJ+BCxeboSyRLNeRFZLEV03TYpjqy
Z1L4imDs9wto7NWVFc7l82Uhp8fiBRMv5xnt971iKSg5k2+cofNINr3BOxi+Azm3Y92AJUTv5lbI
MZIgChxZHnaN9mgiPy/wVuI574umXZCmebt7fXBOsdES7UJuvsCtjbW1fufszJgIboO/+cF8ZsNc
fRvBRlsWL4De4/SlQE0QC8Cig2Qd6s27KmIdT7EOLmXI89RJybCuRx6PpbaTCNLBO3muXtV56nNy
O/SW6VOeyR6u8p4dhk4doleETmheOyJaJWWShhvEE9G9RIzVaSEkzQTXOKIxnZ0mvB3rATZJbx8Z
T9wOr7+MnL0r6gzE09zisFHWaeHSBIGeVq80C0//zCajw4NuPlKTqGZ4fajZ9YP9gW35eEVTkWuE
/aI+M76kj2eFPTcMG+GFdM0OS/z/2LHet2HiADk/POjveloiMGT90fSVJTTe++c3Mm63F/fKJ5XN
kwObK0OCwVKTDrpkPPcke/XDQ0G9It9w+R/qkyfKpBP2rqDw1QWuxZg1JH2SKMW/gSJqppnYb/og
1e8CbJLq3umU0OCWTCBphmJwF8Jw1u7gBPQMv1WnCYPKmeBur15Vvsm2IpaLXDvqs5Xc1D32W0w2
BsdNPtLs0q6SzQKezXRSLvOYhoaFbmuG31b7JFulGCLgHphOFs+gR1AqJcpVzcgafam8V5hdfAlx
G52GXF4hoS8D6EdTzf2bc8h4jnVrlRa+0e432h83L/gXKyAo4EHcmO3UAPu53chCZz8ZEe4tYblv
SNC8JeNG4ogdiXb1uKOV5rocK4XIfx478mJ7mOgaOl7WbLOhWZXBB/ZKFBV1TbGGV11r6j7/66o3
mgKdHxWzm/GLsnqxpY8Zmz/mwpY21ByhWr4KZ8AFHwS3G52kkHBqXe/mFKckv9GXOC05e4mx2K9g
3CPNRfrx+Py3oemT2cVKnKt+kqufDrquXMKMfUa4jl3DoUGL8XUMw1agQKcnKszYV3FRNM7BbdRO
N51loXomBju6VNpo0n4cT6GlJDPcrRDh3PkYu5cyKQcg5DeQ+1/ADgfUUtkyvcfXUNRWVI/lS0xG
wtJRblz30E7Vztb0KG6m/7RIwQUBsx9VGqaehiJRLbc9+A8xTzn6/0k8KzYoDCHS7YYCxywH3hZw
rLxAehdfBHWobmkWpIfIhuW8D7OhAv0/OeqCmAE0ekLYey1sCWIxh3maf78GJr3faErwgSc/RoeB
GphT/1OvjKj34kHy1/b+xotJsAGHM9RY58uUOALWvRsc/5BAjWE4Z+NwrRB+gP4zDfyrm99wWXpG
XYyymk2S1e9Usj/ztuf9ZpzenE7C/5F1nQpKI8015IQ8Sb9u9FPNM5hmQwwbE1QTOxVyTtoBgYqC
BU0kG5nynNDgwRJ/ZzvmeaD0aAuR33/TVxOLrHesQpn7FhIBAiFv24VbqwbOW61Fg+NlkpeE3Ik6
A1ZhhbHSqR067N/4mO61T0mJGo4Ld0ikWS9hs8JZsmhQXiiCjuKdMiw+nfWS1jWPftPECtQRCUfL
L7CTvCTPzCK0kaZh2CKCkMURieaK6PCc/NVTGLR4fU8dLgWTPbAw9hK3ma7f2/yQlmHCx7ZRDmhK
9QrbdZHVzrmnXfIZ33Pr47GEPom4QDDt3pHP0bzKiQa4wj8WIIHb1J/ZjPVX/jVX1X43s5fQtUk0
sSC1/Ywh62hajzc8Psgot/gO0Z9uhRbhGiYjXDg6aA8H6sJOpgYqUun5vpIh26Xj/apUdZXqTWza
5zUYoBuGHbdRqDBUlc8EdScgoN5MRWFLbx9rum+7fwluQmgtYMHaFIH7ImYOfCCGGi4fffvqXqSA
mZFOdSO/njxH3/LMYrhthwe2nyQbz+x+EN6Lcyfv69LhuTOHxKo2Opcl7LviJm8tXUDji6jx43oi
+QvM6XO277+3DkcnP1ciujY1OM7J8Z2m8S470EshEQi1OQT2LTWYcNXSCBI9J81T0sf3VkrWxM2W
gwPHEQo3Tk7hhh7l+0WPOsFeSpGrT7vPhRPVbCp1Z0XWUOk6fQWl9VYyf1QI8EtbxVs9dwYMRd7c
LMWqHKyDc3/7kM9LqNmsINcuQNHsCgDeX6x/9LGoyuCNazwrLDmi8iffR7k6Y0Xu5qxIV5TXHNY7
ZKf79XPXMwAVEzCUUg9y4x4trQ1dnC+TZtq24vJfbrwwPdYxr5KeIak+HkbyVjlVqhSUdI1BlhZ1
9p8zEWR+EplfVdmkL2zvZE9X5gh7Vk4eVIL7vYzTq9atwbTgvmuH8gsMvD4xKIxZn64Be2mK8Efv
TQ3w2REnaWB2qDzEEnDCz9xntpD/VGBXF0VL/rSwppu7mHZbUTsqIsUgf5c8j11TArFVHNJU5uZY
wL86hy+6mNG9IWhtYt1s3/Jb4rxSv7SfEQfWLVrKry0bzHMOFrjp2xS8lbI1L37LzyJE2T/kDn8B
97f7RLcY1LPzWCDTYh6ZasEspwYeNMql/Fz8WM+SN+bHL1DmurlwcFVHVRwoH1XmFgNXLqmcXfEe
k+1ztHvQRIDjlvQPl1H+S5Utmkz8WnrNX7CX+MiS5snARnzVx9dwOwFmQOstWrwpVAeeVkZrTPJ9
aDo9LfXgl/EXgZlfxbylo7e9DWXiBcgrz5MeiIxplqpON+4d3I5FPH5BZCgNRA3c9375yvj2FutF
BkhXtgp3g6jO+8lTS5m+rd/4zww0aM/yliya/wt61WY/3ayvb6quJzloTmih0F8AY4ZPGSpYX3zg
ETHE2h3CeqknwBB+Ev7IJ4a9oxeKNiwZvfox1Ot8t3owbnE+EtVv9jLQ7JFQrG/lp2LlqjGgQHpL
Ng6cnaPbKAk6rJGyopIl3KpBScJtIkMMwQkfK0SBF4ePEtNlh9OCkLkllk5liaxpXQnrZ7zJwD1q
6+6wLGKXksfEN6gS3lgsEHCqkv0hlPtx1P+an2PSHUozDUKb5m0Yh/h12elq5+z01Vlax1QScawc
dvtmPygKIuiRsfL+BHaIFL4LFlmGf6Tl7cMmaAkSF0ZnpUynze1Jv15LPAYidoGErjk1jWZ9w3If
mBIqfUGGrqn+wiimzsmQSqLL21l1cG0eyZuGcbfOE5U0jVKQIn3SjgKlneNrsjEbZ2Pqk3L3DZjm
AhAgQGbO5I49itGkryrH/5TKRhjIp8+ULHMg0tY1rxNrG3fnfFvpix/CHq6zjDaKIQhlAJJRqn68
lrTLJMUNDfAexdupie3cSTPQIP1rmlYQY+Od+3ueKes3Co7vYUlF7QcgYveryk4+2Neako0OQSl/
6UTvXgHzH41RxnC2RYgzIZ+aJHAzFPaQlKbnhK5lEGJiWvMcNlEYIxm8grnNxIlshMPmWaB98TZd
hm8eArtYcgMkfOpDkBad3rWnVyiwP6+Hy1RviDRwCOtfWjs1h6ZxT4RPs13PIdivgVj5Nn1NyWkf
Irk9jOysvZEU45Q7kAFqCd6NRPJ1r23DQHXD4ctrTZYzHKTKld0CvcOJnBUeul14uHXhMNC+EjGv
qfKK7UzVEcbFr2IEFMQQ+0YYFsiBkNropJvnUX/2pYsgYXYEW5FkHwQOaMi2/qNSfrPfctqitHUq
yMALp7TV23hXBkE0lfgZWatCskOIm2qtc4GXxDJ88nuh1I8LJbQRQb8xgjVnt+7RX8xR8KWLEBUV
Uducu6fSkcof5cdefm/D3DIXboHOTTSiz/Xtx/s8JRmZ2H9gFm0I9ibEBOzJNXIWKfqRjwto9ORZ
g8Z5IXsLnrbJzBxUYipXDBLeQAjJxx9JZ4LGd3ld3F7faJD4SyI4VE8hwt/JTCH5liMBO+tM+hca
uAva9YK1Y93ySg6jcZ/b7XqMdDivfO33Xtw5UHxyI6E+7PpKjwJ0rUv3Npt1WhbyttVv31DVeiz3
VVwS6f8L+ZSoFtWrlBN0BYlnDnCE1150QAFzS7v7GRia600OAoFvt5cxbCDI4t4nGX88wAcSa425
Us4QY276OX82bC2xF1yjIVs3LxuVCDDUwySIN8J7G8mWynwXY7Ou1XbiUAS2ePtcVao5eU37UPiD
+iPeHfSSX85kur93m3f2372XvZ5tw3vHjkzlURUYrdDENqD0fGRx0s/yuHBZmdbRYKifTDeWfA7Z
QoKODwO1gbpwFX3EfZGmYUldlKRg73Uft1kKEGdfJU0JpPnFzehq8LfoCH6Eer8pRuCKnpyQteeD
nLLH6VDieExWb5cKrP1ZuLRmlo1NASXLYipKxVBeEltYyFzCAoVPcuZdx+Z+1WVW509wEiVj6ILU
RnJlPAJFjaJ5euHT61VyodsFwIJUYLSJtvfQBswYufe6+4cs0/hMzRuvPw3GMsecmx5SmSaLK6eS
xEF8ujDEnkcBYD7usxY3Y5ugxJUdv1ASpug2KBPGXySTvnt2yIY9TPzDqyEh9m0g26zAn6s4YXMl
HoIZ+z3/F1w4S7yNicQtKnZOlkIMSuH6biT26+zlk2JffTAFyMwG2jQOPHf+N6p52d3mi65En22c
wfGJTiyXLDAZIgL9132Ue1gKNM/CFVXLrLAdMERjbrBzdLDPqZV2MMzUqM2ftkhr8QZjQ1r60Yf9
RJizFCeXCf+rJmT54imVM4537ELePODp3FCHEIEAkVyLMByAZYV3ydc3DtOBop1pmINOPeKBBBv2
+zl0x+xTRbRE7x1Da8j9q/hzDCzUpH8uB2MbIpQXiaLwm6CauQ7dD7ZqkJhTN5uX02uELJpTszkW
wvXjXRc1kY4Qcg6Kbg/j1PTGWlWm/BSsQst/XbHz45VJd6t6JFP6yU7F6Ni3O2JQljnwMnebemJ7
E9syLYIzw97OQr4XOkitoIz5i8OYlhsZWkp8D2owk/64t59F/eDGKSDaiDvT8yeYElBDOP7r4g+T
qmV1gRzloexQMWZaD45INkHjIRXUYD4RObaof+GTHMoZCkOKD8abpPLZkJ8Vnn8zxVGiBgZs4eKR
E2Wn+6bqkV8B1uBONO0mAZFAyqHBaLgvf07SSoxmTOKXXQgHG14ERTVbJgPQGTdr+0ISY4SdCbYm
ZV6bsbt+84p6Iy87fLA4MFl16PG/nAssRmdVQw2MwXLbQKVL/W94TwHqo6ihv7xSSkN0d1mdh2Lu
EgEAJ1C5tKr6IKvLcwcMk4loemshyCL/Km4krIrF1SzD1aT9uFdbYEbm5xCVdrRHDDJJXoxP+k7N
s6bB/pagvVkmXG4hq+uT4nKl11PiTLTIA/JPQ0MejjIk3KgdNWkLh6mGaQtvMIPHiQZThma6QbRC
dxU2GwMGDAWRgWN/o4h1L+tOEP7BhWUDRRWZblRq7fsWtlXB6jGOpOMHK6juGFU7HLVWKPZKloOe
1KkJgEo2brZqjPCsS2JzPC63zf34PvLnWtOPgTvOIx77srTbhQhSTwEZWnaSKBb9vKEyl4c8ruGf
Cy/B1nzWH6FTkrskW7bwFJvh8GUzMFKk5P6izhnFIVrZPjHWY6ZQ6PVB8DrwvLTRY+5ccfuPnMbX
aDhFe4VeB4vJgEa7VPktdHC71MSid/8XsETO97pQ9Xy/ba9hKuBkvw9FPBGaC/LPGvzKjjeaL28u
n3OMWgefwJLJyXqwYuSeVcky11f/0oHnXqwJddiPwfhNCUuf7Mg7I98YKfRn6tzBh2giTLg4eCNv
3oDf+gWRgB+O3DJzsKE3kx1s7e9T1MTa69tMA5ZAXwMfxxeessw5NBqWV6JIDv54w2Qs3z7mK76b
TIveNCYvw0QchyKt+fHXQrDun09YpeW9L5/cyj5VGYRx+eiF22e87jr8dLwwTdmtM/fkQs+02pty
mZxnz8ICAg8iPjsTTd9BjQHztDyudo2Wa5AsTkA6dCzH+bxbUJAv26RQ/doMTcAdn8fIIz2q9Zr4
KlMDiWIS3bYju2twhN7ulb/RtjZXdeaedYCDEAhOdRVsL+wwBeaT/yxl3VLUISlAX1ETf4E5cMGo
HS3DibCo8hWGx/M/y9s9K3NicwYWFiBsjGcmmUXM1WTls52CE6DX0zPWN/ldTUERZSOXP6mIjX1R
i3lvACUXxrZvYTTnhgKf9OrWRFYBv8XSuXvNiEARu106gBH50MMSC3phwhgT43CNxwqnZXBnzTzV
K/53zwMuk03T7FGdtvssdXx/c6ZBfdsBdJeBlz+bP47i2wfNrzGL95rG+PYOMxj/eOwu1HimHUhX
rJJX/sFWtF9G2ndrKb7lhcHaS1icuQhrbAyP67gKAJYb3SHDE1TtyKPjPRJn1LC8cu5zpSdZ/jRr
fGFVsBvBvr6My4URewCuaxeL4hT5LtSxA1LECTEacUft0mGlj/0PuhfZ4KG7WreZag7RpRczKUaH
Bj18V+yaMg9uJjj7w7Ec6cAbU1bi1XL5ErNSW1WzeftMLtRKbI0YKKevSFGZ/ogy7tKMik7KGDhp
E+LLTzlcYNp/9CLhwNhHwd8SQJajjndkF9hs9zSvv5jsW5hvNFiqFVPPE+o5NOzkXHw/s230p1Gw
XWf7Put+nE/O7Msix0/BSu95uMU24D0TQITiMfsD7UFdxSraAAAopfXHMyPfTaYjUUHGuRjkOrNt
gl1Dx62QIT5mRTOjEeMo02cWsq8uioW0EwSugqHScIXruWFqogR+xLCtOJwv96NbAWnUZ/Zm529c
OHSWFp0n9GznSj4tdAp1szDzgAgKGcELaULb6a/zdrcNYZkto6L6dX3VKEyGAy/WFWNqcQ3SpudD
KJDDwZzPMR1cYWQpqcR9m0HqWZ3H6f2ne5s6dCLvi/AsDqrtcBQtPAXMv0/5qhnBVpt8g/pah5bo
chN7OeqoaYNGYz/89iGlcT9SlCR77oeWv3r2PclXrBum3dPeG5g28suTO0OOov2ofPATYaDt28tI
qIMRyUnWDHoNQISpHodyDjKbYKYnxCq4QQdL/QwmB4QQOPiy72Fgl/iS8jW97smUIL7ds/h+wtZQ
kcRBnR9L617XqeTQ1Xo6fjBgJYEWorFmtJb7v1sLd+wvMjnTPpJI6+9INEETf2v6erbV/bcl5RU/
WOkByjllqSoUj9w+FDGwY7k00uabowO3X7ExSTq+tk8PSDLbkDW8E6oyTYP1Oa4HaB37PRiA2v0t
QXmQJuPva/T1ZDdjHqk7+aMXkkexJtANWnMvWixO74LRRJzrFY+x3rUKrclvNmKriKJms+hjHqQo
ci/oNAJruH0K9G90M3rH0yFNVmBJpK8CUn0yktNTpK1F+MDXNPoEYQkgrPROvvX2JMdrU7lsWpKF
btmQQqZRyZ8d8XENlJKHJUq2zSGs2caMLYNgtRb6fXHoKRyGhB0dYhX+KlY2tvxoVoVffP7gbd6N
BJckpc6dWc5lHRL3etlWa3DQjrdQ6/WctQEXT2X/KNZZK3Zc3Np5C1ZqITjybeJrJZZrSqjH3FGP
DXWX6W1TnzkzvPIxz2FqFi0lnSEdI+tyBjV6M2ov68BCtoNm8eQ0KaFZhCiX0PA95M+x69W55vfG
5dLeLNtW+gWmM4YfKxvCJEOsjC6gQp5sWo+jVMWcAR9wRZjWJOXo/S/9+9MPEvH0d2csUQHgzEK7
rdVvnMpXjw/L6TENt91Uw+y6rM6+y6IRlcg6HafPAjNMKkDL4vuXaGacimaxG3Z0qOHlkuFdyaQ+
6lF/+9qys5adZf+EVTHvXmRZAZGGACNMkxoBd2CJSlBnqmG2BFVOU4FFqqkTK94fXo6AOsyh3jJZ
TkLaSIxmws7MUAS+Bq6EBJuWhno9ferfm8/b0MriU60+T4F5lAXLdARCJ/SOKC8McovDuVXis6+s
xo3jkxK6POEK6nDPX8dFMXyI+QX7CpK9oq3w0BhghSrm8yg/8STlTa7hIR/Sv8GkWInxSDLV9wI1
eDYQ6iCFriN7jwS+Ipm4L+9A5jeNWND9OVv+uf+vEkXPf9FOuffcAVNOyWsMq3txyJZE7ZRt6Ml5
L8fayw7dStKrnsXC621IKa/VNbgOLrAlmgLWtjpWCgEt/aHzRSiUjApZf3JF9Mx6ecv8lUN1vXpf
OId16E+KaGrDEjbx77jzoPVQOJH/SLf43R2cSyyj0Fhc2L6RJiPKFtBe8S6YRKsrHWdXWE6jhxk9
DSLcq7HRGHPRm8FTfT3fxshHFK25bpsM6m7qkoEwBEB7f18wayV2ejXdxv+bPgyMMhBKSj6LvXc6
3dCFCk2xj8EARyHaIS58s4g9n4GeI/lmaFVLpo8H1WawiBYdIoWMFo+DmrQ7EV70a1i32SaZQ1mk
yqf3c5DuCxggXqRaaYtOiRAleYQuxzLutuh1m7cTDRyBmduQ/yTVD7K9Z5nZpvne0heKPDm9FDQU
TmZwVyFv69pqGVA8MbhYkpHk1+KxTOu51s9470Q07Yn98UbuadD6/j46XUjGiGBcfYtEochlPtGa
zJvTjbL/B0Am3bl2298TwbSlr4jwAnY6kcZmU5Ydg9M6/Mtvxc7f10YK1XRoJ2sWIQKvicHETSgy
qGJBwj7Hr4fSkYU+DS44w2by1uCbGL+VB4RMAOkFXN2yBC4hx0Cy7XUzLz0KdewcE/LSBh4jnwf3
5GX0etAkYpTpjhIH9Bsqf7Ugw9jbI5NlFTFcn/AKVfpvzEfjEUruSVyvGJb5G54rpuRgOlinsOCU
yam0Rv4oIPK5VJ8jCvy0dxaOqohOENqrSpQg+wW8f5jKxHn7Hkcva5CwJkJN6yhdOgtViMC3BZ9G
Mw2JeeipF4kxItGU8oKly34fpmTPJCN10VThVdUF/BxKOH9xt2b3+ic/bSIAc9gKZE7TOccAyqei
lXnUnTIvTWe095SNDMVsM3xAiKBs/FWdgoRHwdi/PUQpYp5cn4XQV9ZzDVPLafc6p3DwZcyVtmgK
wqs+yxkTQ7jBRLRGCWBpfJikY8EOzRG5uCeLIqaH6DxezUWh4ojnB13RIKYcAefYbs10KNPb74ND
0325oG/iA6UM/N4wbmn3YDwV0TGTHOS+7QJiV5ebMdfFGVZGlm1DefVsJ+eoMoYvoO4KrXcQcvwl
U2tsm1YSuXftHS64CGdIJPNIXFMOmNTdFNz7xEfknqgBAYK4iHnyL2+M9791jEg2toGWPHvXIkOf
1u/6ss0XrwLMkcYbXzCIAVHSsGZOQDbgGcvDavmdRg3f851p5xvxPOYluhi/5+A2ERgl3KkyftOi
wtv6kUQWHaRXDO11KrJjXw61Q69VpuXVDiko7zm5gjZXbWFra4YvIdOIO48/GR+CCyQVkKSGfcn0
IfhKlERuJjDG2hoLFjif9MVSUKYXwEwc1pKNA0JdLxspufG8z5zGyl8UgplCBwfSsBG0Te9kl8n9
EqQahRQa7P5QnrJ4SBdehxD1qFBNTkLb/pxNkdYnOJV5HiUpXyGc/JKQZomRAB1N8w8MAw+n5VMQ
oo57KtNeFSrKZOPG755i5x2sx718V2SHJM9/MYwLqTHckfIvIACundylQK/NQQf5tpmeEyP5njpA
MXRJQC/3eC3LhtCE6mr4W1LIzp8lu3TbV4TEeeuDxrzYAwIvFkqwgBHnbDaTObKcwNMcEPg6nd5R
IPvku7QKEGQ37MHk5ksPcViGRnqw7mASoYyYquOY4R6mPT9XEdatRDQDsJSVmqq4ZtTRpzluJTvF
vD286ZwllIm0aEu6U6PVBVkH9UkGed8o+LJKE2fGiabmV5SV/08fve4BG/Ba2IA/TkCAxPOSEOMb
RwfJRB02GWxb61CgCayHmgjnriJla7dVdLP44Me0+6fuBrGKXWY7cE3fFoXr8re2W+67qKvA3LEn
702JQR73VEuwagvOsOeu1Q4r+JSsZQ+9NKlZaYykzqBw2kkoRQrAHbyPWOB3mmdjdyWVG64/eW9m
6tPUocf6yXXKWd6uwKU0KxteK3G7q3YNItDATg7xssgs2KXUTk4B99qrwAOjnNfcESCg+0zX2b+6
z4Lq3TjsNvkH4G6Yqd6+ZMRhQa51NqUeLukoXzxHC5j0VqSiVRWIDG8jnX08Bx0qQhdz7Uulflo3
9JK0TZXhXkv/yFBXWG9S2IBWrJ/WuGuYYxJKrvzD1Dl67uUFinRLnMDmI3jMTgKlmLxIxkGgE0qL
dRVqg/HIUODsrgA7zd11/p0qE3QL2D/alaUm/kWXk/cCObYTchxX1pQ6AYiWdWbhsAPQccztVO2i
YceDavyzKnTD5KhPnsRJ9U97UD9XxCpTFPBTGh5+h4yXUv4KFT8R/tOKiPv8rBB95Sp0ULC7fvOv
yXY9fIbZMot1XHVAsLk6S1hT0dWj/N75AWgre12QUTw42PyCaBFwCGO9suMgIakRhewR8kTYZiBy
EibPKiVKcTLnP/3/P2zFao10L98lBew8Ck7Orx9CnMXlHnMbcpIgCzEzqGP8oZNGIzv8FhCTTWPK
MgTFfbn1z8qzmgWkO7k/KGdbNjorB4B1RQy1WZu+wDGv5SiD79o9h4mY/P1cKCUC+V8II0thfwjH
0fFbZxyDBjdRubkEj7Gpnw+SLLlUVR5RB2jeAmfKsYu4KhO7yi0+LThdEMEaX6+s4oNG35IvJgTB
h8SJZz4o4J/4ITXkNaQl7MkyuK1uLEOd3BfV+8W0kHsgdZDtN6u0hoLHbGz1ZfM4NJmAuXcZ2eIJ
N11N2sjHR9RA6r1zmqxAggaWdU1y5BIsEXm/oXRTqv6PDyZj0PRHploE0o4CeukHqv1+tK+fDyQV
4VMJQrwuTydhtsJZH4maiIx5C0fyC/aSIbEFG7OLv7QW4K7VVEKbW7jNo0NKHYnnGTS5stW8XFLA
Q7TbOoYF1Lfc8mhl3BzB4Byb/0blKS9iXuZk8WuNwM45mIIPreTVokLVWmTeP83TF0RV5fZxEVvV
cnlvmUsLiI8kokSQYJxQgwjhFOfCC/77Es0nCn/ezo3Zvw1MXgd2X4glddRISpK+9su8HMpANcQ8
8eu/wt8odioOFuitMiJlKXmE8efmlL3caqflrLkXedgCv4U1zEkty/8yMJMqUK9O1HkZPkxgDXEA
5FtCIZlbf2Jbh6m7LYC7i5YjqZojyqsgJfRqr82RRCFbEvbPJOoNGaIFDP3pQZ4sLHPqZo7FYHiu
JTHOEZXTaHGjNIZb2iCgra4wh1frRYIy22D8zv1UvUZ0aUcHz1QgdetW7Rekrx6qs9ApNSukf91u
/GLqYnx1QZURf0XWeI753J6lEbhSM80kNThS+u4eNtWBVdaXKSG0GUeo4VQtbWaUdGcoT77s0khT
0A6sbIyMUPSCHqpLwRF2eKYVupgFK/WtRDxFzemGQIR66PYRFMoMw8c9SIeQOkgrbKBTH5XzhkBG
KGHlVLOCtNHSfmKVHbHuUgjQMgcptXDgu6nMfrjFter0cjog9DAg7iS8zIR+tsGPWXNt4jUdq33Q
hpEv7ZJQ433LcsvwoR29YWjkZ/Cx1fSw998kie5qjlWOFqTVxnXz++QHF9zU+CdW648LoMxs9j+A
q/WzBc5oQu4bt+PX6ysz4JCx8E+2NhC8WLccTBqDmdslyM9c6IH9SDvaYK4u9bBfrzoK/7SzX9qO
/3YOXRZ2GOtinHGE8V3MLrxaBD0EGZHZDKjkJCrEP67VzAfT1YrZ1Y6YJCCR7KX2iWC1rnuuvlDd
7OkN/n8xQBF+0CGki39gbETmKWjaC2wvoBVKr0lxbIG5Qfyt/+W33VJU/i9DpDfUlBtxxJbqgJ59
g7vwcWES41dWWReC/TdhcM2CzBfQOXbysX6MPeF1l1P9tDdS+ShJyr+sUVtI8MKslCKFp8QLJ3YE
vp8aH5vmNMYz4EvzAPP770iDmgy9f8dHNNDfwAAKMFoAkLKtUgebidQjv1nLNJyoQsDRyqxJ9Idx
5kva1SMXpZtcTtq1JeyyWDmHqFb2ecFxMDdnLIq9DWXqMNJipBU8YBPu5DrqfGcVYq/mKZPhIumG
UCHjZMy2wULU8GGlHlKtXFvxWhaeuWOMxy+rS0kOV0KAFzucUnLgPSVd9AVJKayfwuFKw6zf3hl1
ZGuL+h+G6noeJOM+2l63YO7Np/vjc9rHxnv3NkqWXoGSAigoH+6YU5k+SwDIUmPZY/7bZAI7+1zO
T/U2te7Szk1rQeHFEarZUtooSDEyAULP5m5kluCeWcUMDv3eLgrNv5NzYPAbQeHLR06H/vvHYbS9
WYC2rUasapIae4kxlsS+2w707Oi3hGoj6EqflHlhfUbblYG9pZ/zgc8YuAimLRkUDiOR7zr7gdZQ
tt2mNVnlabn8am3d65j2XfZ3wqkuTIozIrl9uxJTBtT9X00q3ClSwKNxmbo7+GigjfFYfsKXnLqx
euOLIFSrq1QuNZJVdghM7ioK96k6mJJ49G2A/XNFhtxR9YoOnCg1qSGaiZWi3jnGQqrYtj4EQwWz
LIgN0iw14T26uC9HMCJCLuye63didPPWHKdOhVU7ExOru5aQ/BmGYcGNelgQ6+zb/2SHtYRhwnTC
TJGzOymdrM4VneysISHCmUgHnuDYJCq8d6v/4RrImo7BIu4jibvcb1svSSsQ6DE8TCACuTRTLikj
7fbrWPMMwkTJ37+8a5zGl6YWcjPfYpEjF19IwoaCsB8ZIlbr0f9M/aiFTGLg9igrfHczxixK2Nef
DBUufIMhrKcSLcpj9WvX4Nl5PpYMHVIRKYQzn1HmMJEv4nMPREzcn1Y2BIBjh1ZvT3uUc4Rmpm3G
+vn90HSb8QzVNi34TOiwV/wcTWuW+S2e6HnSNK0klswmySdpK34jii12kizPeFOfjsbhLrAMnv1d
tNdTctP6OmHPywGnJ/0X93n0Z5VCX9oI4nk0tgqg5FVBR5xFXeL38kHIkFonImiJSucqZ+KKDomM
XKVvHJxtbu7ZbVsUkPkUnMXPmkRCZadosmShtCiuPHZxhiftt+xTd/T32c23uxjagIsq9O/TyHbV
KeiLeTYRBvMoiBsfXNzRbD5uMs6dA/vjio5QP5QDTTDWDJH1p2IW5w4AbpnTVmsrmG6H1e5XerSJ
285F/JjmdUcSkbeuOwXlbCspyLzLiWEoR3NNvJlCHXXHnW00hulrIGcQfrqzoeJm9I291555uFo/
xDmSNX+SkOE1dUBAOsO+5htPQ27M95wJWZtFTyy0UN0HAR9RGIfmUeGLu0nlDDsMGNlqWviyX01i
vjQa6pA1jdl3JK4qpbImSZ6G7XK06hiRg0qJEFrOpgkWcc+iH1A2t9y+YcXGCIEKFkDRAK779iUe
dk3xle0/GQih3mRW311Bf2kmtXgdM1nUh8Grd5qDg8fnfaAjI2DOfCfu+TZwmKP0pJVkyvR5VJvM
Szvrp1k+KGaIJ/uYig9YN1OvVG9jMZ9VBpM/CMaH6oE/lpm4frk2zGWnPrZse8Mypa17hU4wpxNb
lClUXmb6XjGINocE20lJcb7nOmKuLm61zy/EW+CzpG5oqga3+O82Ar1IpUpdRy1gMaWFBdyS7SLe
6jgEswD/jsKSpVcg/skSG5QHQXvzGJGEeJ9D0u1Y0Jf6YvLsvIdBYof7Tb23WfcR0VAPdVyjGywj
MyV9tgUZiXIX2dLp5d3Gq7yToZaWeJuDWLGs+GR7ColxmasTM56Waj8AwDJRLUM/Y8yc2KH7ow7y
8kYR7Phf1eKV1ctaOQPRDIfgc6L6QHdHdnP8P6Px+rZ69qdMyLvuPJX/+zsFiFxvvZpmizLGPUL+
y8DGng+sGkg4Q0cS5XZnSagGPHkF4K0+kS1MVkz7+UaUDY2FGAKo2S3AtMtkLy4Kupk9VDwfArrY
+Ma4E4/pdHBRFXnO02K0lkdUdP/KKU62joCxd/ztH95zt2eL/hR+nSo8EvJjVFAQDAAKadOPBGPw
FmiG648HQn8k0ycukN52XYVsLWKVcVjmHiWErKU2idU0J1xTsdHnu4LbdZ7vEcuaPWDdXhlr4vq2
wt/8eu6A+K7A580LnIH4+Us1YQ9Dd2S2KolW5/+65qY5JximrAJw8mVmlbF0CwjfRvWkbZX1KiDa
/rh/ZdiptVoN+xO8EfMYdu+c5DHN+m6ecKQqboImxCLQIXvgyzuv0dHgKUXCsqpglZXpn7KVFkEg
3YgwCoHyvGzGKeLN3riI+Ve69DUbijuZE+xq4t2iKppe5Hvl8CxnTKK7bdZ0Gjvl9HQfgFzkODj4
NkppD0ak7xHxdKQ5GRvn8XbStOMqz0/ryUrqS3dcNaxJQzvEDvIDGV9vNySKrYzzQR6lBvUkVqty
sjVVGBVb3GyjeBPudJwG3eIqMsLZWqjVYe/t1w6Y6yaRBB1cBQGky1WIKMTqok55nfZyp1dcT2xA
iT58+6PqAEZtcZFfnl48lsjy0OxzNt1rwXuPDsY14see5tDTmgo0NOcaUWXzclkbARrIfMUpuiIW
+CaFcW7YbdfADRQdE4grtgHWyBfEic21af9P15M39o5eM2bTo5H6ZXeuaWSZ4100Dc2ko+/AHR0a
FHMv5kc6mgoAkDa8Cilu2/GDKbv/VodaUYQwNOl9yjQC1ffIfYp5zXgYJj3oGi4ZAdQT27fLSQnv
1arQiUN7yuNSoIDEmtKYl4mIYVvsLPN7V0SuMI7YQp4ac9+BR4bVluCB3H1pP3mOvxpHQ1EdjS8i
4jKzeViEcOQU+Tdkhx2yOXzGysu20TIKDptrqs3K7KEHvOXTh0OlsYPqxrxou6aKaEq5gfbl34/f
7zBM4jtO7eHku8rrDyJw9iPe+c3gBCRO9iYCkL2tWc6F+o5wVb4Y2vH5/r0OhGCUUPQwCBhMDQGm
zWCBROShBNVExlIM9kgjz1tZrgyC9P8ZVl0koaPrc9arrfzeCWidhagPGxUQebGyLLBpyRteCE+9
TjX8k6ZNTOGLTCgG4hs+Ta2LLSnd9tZlEcf7sSEn0sBqoc+QkJRIaN5eGLFRVOjpWi9FydbRF6D7
6C1or7qBcxQk2R3rT0u1+mNkspgUe2bKuHH+6vWc6tKXvd95yBMp/TYM1hxhqmpnVQQnA23y8Isf
BkzekW1wJ60o9SGbbqnhnXlM8FV6uOJZod+0e/wNNVD+bNPonFLRnXuXUkiuHs2xaNXBeEIiwv/9
lUC7S/dmVA3uWtzDRStgMiVfa/f6cV4ttabg4g3FnYLkVoVZyyB01Y+XNpSLK+W3RDWYeOBP+WsZ
sPatujXCFK2JDfIB/mmJUpJ2L2fPHIHfhJGOIeAXgbVySx0sXktY1hocPOGl3Yc/uGRq4rTsPb6H
s210rhBslIX5rEEXns1Mctm8wt1G9DW5DE6sBpySfK3jDcXm/J9PuPRDlXoj/CkELBB/6f3JYY0U
hegNMsGzduh8I7Zo1l3ou1YoSaEEcXJSYzX34Vzkjz5RtDoPMY33AiaPQ+6czh5WOgNIv0tKhEpX
2MopxAi6W9g/T+Jizp1hR7+rjx8JMeQpmOxtotdSPa/1rSPPC8km2y/ODuR3D9YkQoYJCw//xouk
6L+pONZN/bQJ5NpDz5nyiAKd8CesX2JBXJRZDGsgtuUCU2BqJzklrPBWYwdFLXkTQIvFrwKGh9gu
87mvPZuIeUfgsgR7BhdzTIShp7qefU+taUagive7hd0nCSGdkneB+xvB7FnUmv+jkpxM6Ug0oC3d
dPfzM27sgwEAJD55Oeio8QIKFzoGeSPtWxgZwErXXFpd+8st7ajeAzkiIy8lDT10HPBaB+OpdGAx
Q3eyA0uWmr950xcNvUZ/nbp+UnYTlybKS9TeaoySKPn1eRqqsjOCq82Ywfavq7EYRqn9Oixn3fHs
9NJcNyzmA697JET6vxapUrqoceL+B9smVGDb3OdFeKwufrqYkGJ+yTsvGw7IuW4+23ScqaS+Sbbk
zlc0t0EjcD5JCse5caW05u4KRTyC8Wkt8Hf4eP4X+N2anL6jN1gZefMV8IcnRDLqoitqhasXlyUv
zPRPiXSAlThEZK2RKnsAWH0Lzavg9HZ0W53q8BRT4GSyVSxk2j6W0tZBeY9wLE0rCdO4As/szolb
0DFzjb41Ik8RjTGk9jx+OC7cpjQWSEUZJBgNuTl7GlYEMxwsSgntKLrK0CTymh546FJYShBlsplX
PWpjatJSEnPxk3fThR3yfwBHR6MOo2so9vZjnzTe+an6Y57aGzrUgIEcivdV7yKh7UOySCE0CB/d
UkEt/qIaSz28j/cLqhMWkYn7nkARo7NEJYQxIZPTcRo9ApXK7JNUf8XHKPCb+/M9mJgBZpsl6LRC
5evPm86Z515wIhKLPGToYB3b0rewUJCFDucHBXAKJMBuLEcv50S3Sym3DYo2W3/4clMeTlVdRlod
J5X8MOzS3NrAc9zfOsKsdX74WuFsdMgFMJMgUYhx6z6FroTfrEcnKWWGqtgZNoKqxuPffpu+HsNk
D6Hqz6B2utZuQG9bgEixwD1u/SaWl5VWfo8AsaRp49h/kkSt2aivsaAoqbwLxvP8BHTkOzs8X97v
MEwFeR9u4QiWL3Dgh7T/gGt6q3jBm4qiHdDyDsKCh6o7zU0BLGhZ0pNVMS16riaOs0U+KHYdXSHw
xSoG5S4qwo1nvIC5HCBjty/E1mCPagSE5iOTXd8z0JrbVtFkLJjPpcnNiuCCoiF4NlDGciM2oTQJ
1J91yjT7emQNmPD0PwOKsUlm7qjaAqMeYzlkuxfvVMamUca8oiceZcUYvhatEDbWJp1DqTcE5Mwm
Wa/I3phEZa2fvCruBkjaL+Qsd1l/OZeO++lOSy7M/QVTKG7hcmVl6g0ksDhBrDJ6xup5roVVDmzQ
egd9SLHVhc8ftew4KB6fjIDdIJT/sDAJKkohoox5Vkt8wli1wc+WtqD+ixNfiu381fm7nrWlc3nH
1LqpiCwmcxYVz1mahlRgIftJbyYP+Nx+BIo0HSZUIr5jtIqZug+3NRf1Ebo7lk7KtLlzmXB3ai2P
vX3w1X1KnOfwSHbTvlTj8GUZBHezO3WBIuhaVNMgIOreRlGhcfk13iq/42WJrQke+mnQapPo2DLn
KN1zsN2DP5xYKXE9QVjm2PpJGTeVzCawkaew/HNP3oa3dhlHrvF8D4tG1I2/ESSONa0QovrwP+JA
k7lXC2KEbezmkwglvSnf5HVnEPhiQgg4lvpHeJ5wiCoAfd8EaqrOboh9ghqqTAnFEs6LRzUUKEoK
56qX0He/UrjvmEGSGc6kn+WsoG7GdlRpKKt5uFUbSXdleqFGzijVCtMDHQjgibZRHZHmmz5L5yd2
JAEKjOeYEQeKuWPncdB5jZ2B7gbVhhiXpf2CnAoyD8dIpC3DHS6qgAosA3CGHK2M+R4hbYS1xbeF
EhhDTWl4hwsCPXN6uRCW4tTeiLi5ly+u30RXoeFiCR3fuMoxeS6W2nIyxv6Jd/tlTM+AgBFQVluB
Uk/TlRyWz9A+iHjdWWUF9pVDRYP9dY7jD3gbpoZ8XQt9e753CGTbOf9ZxkuSck5OvqIc+3EmhMQX
NHXLHoUPeFDdTJffMx3VMi5BjE3rfC8ldILazkK/gMV0af74a8zvKSyEMGMdOCvK2Pn45pf6JFlY
GHjR4WBHVKkfhubQUy0XIIxqA4ebd323fEuS4OL+T2bXD2Brdyw2swuqUhTxsNyNXCn0k/YSruzf
9Oi+HO86Y4W8arKS6mR45QneeHVq0AybCGRAcOq6FE+rquVWzA1/K3ZI14x3/t7U6D32VE2TJHSX
ZJmy/e3L6XKkymwcu4L+Xl5az2uCzgSV50Q/Tziz5BFpkyO9+ZLetke8tn3gV4+uorXwVAPtkRXh
7NoIFghwbqGVTU69uP6AkxNIOESDERZZoWfax7bH1G4e9zJYH/DmTvm33m2uP7tZu6Qojk6VbeoM
aoVXQWs8xXs1/gNIZ5rHMgatUMsqoocbqGbJNkzYTRx3tWoE0K1gm5XUKPkymidrqJIOCzlUfduS
+G1R8nCERsS0UEdRM/4qnhswsJchm2FqP/CWZdoLJyo/WFw7oz6ioUnUvvC2eljqNpFfcv3cH8d4
rDcFqOzZeMC5BtKLopYzzv74D/m55tQt6RDZu+9njIz3eV6A1rZxvV5Hqw16VycXkAfStdfavZm3
twgLO7awcViG4Zk9kth9zXCMBvwqyNb9XMmVycRaZkRsDMvL4SoF9SNvE2mYZmGrCEqrV0iU9pUL
lTM298pFQscQizgH3QX4aO/owDPIsibwh1ubZiHuDBzdLYazj4GYdzm4i3vt99MMhJMZjRTI9kit
ra/jCZkTMTsARAK0+MZvTqB4HkMKWvDziTV9EgoCJoxc3wxctq90yF61ovdom168MgtSDe04R3ht
cxy7awEpR5iHiWTlSaIm/Xf7FgO2gUZRjRLIm5eSBZEdldrxEu9Xog+m+SqFcLWCUmj46erRWd1B
5QHF6K3PhwaEt5Qb2XXwtg1AO9NrCUqRfdGP7C6Z7HTPFK24urjdBSJQKvWOcfucb7QdGrqApQFt
MNv9/ap8IUKkdByOykR6zcehw+zXlDroIfTWepSHkKIMdzryNCc/3AbajlC80bdRLlYHkgmxYPbl
NVTs3FcVsU55TAcde0UUBv5H7z+TWvQCDRdt1wLPEcW14yUdYgAOmLvYfeMEj4RurxUGImtJmv6P
VA8LTkF2GioDmf8KV6oK+S4UyRGHYN5pukuy2XZATyEhEme1rCjBCcYXfymyvWTkKFZubxESc5iX
qlRzHQ/Six7KCYUZxCXP61qLuOSMU+upBLFa3ZWFBTcbTF/N0Qsanxz1y/hJNsyNF8rf31v5JzQQ
PgU6k9d8vZFxspUv+7YQyys6JNcimM0cTutLww8w+SnmBGzOcOo9sX6Y8L+MMXskaJ18NTPrKEpW
P9azFXw81D7I+6I7OcpxkSW5/SQS8xGX51aoeY6AiNVcFnf9NC/RpIcb/1NvcyEuZPd82Fy7nwYA
824ihtRC0WXz4KOzFjCXEdaEM69yuz4hiEwk6ZYJpFX91rGspiHwGFXZFwZIaQbFS+TQwrn7DPC1
u/EHVukZnYdx058seKnyKb0KG18xmg4irtrx86JK+24484dFGP0Bivp38N5zV433rxgTO7KWGGad
Hf1KYbS8jJXGoAKq3fXqtXHjnZnWwxoge6pMZC212aNDDw0KsnkI1tDTad5s8WvliZHjXCk6f0jf
d+iHbiWI36L696JYt3z3A/gtY0J3Yf6JYcM0TSlSIifKOD6wlI0piYh4vbixRXSsPbM3aO29WjUL
hgotLVEo2sqcUVVmIuOA6iRsSO7G9N4bhsmQqYQO5ZVkRzHiA69X5Q0ao3cMxDYtiMAfyYv+NBhp
s5tUCbPZoPnasneLoGxwVa8lml0h3YXboRxMYJ6akjr8Mgau6EfV5G55oX9MQ2RXEW7dbj+s3MZN
qFzATMIqHbzwGHvLKT5I8QR4iJ6Mzs1nuqDDEsx1DLl6rP0LH1yAtabMCdP9+uVfiG0rAuQebmWG
SMwdpncgA56QUrbtShULNXRf4++8NQded4T6iliaoE9/XSAaoSqkwKIMyLpT8+wAI23M9aL8pVoQ
MwSGhB2yRgTZY+UPYLAntGLvSrDx14n03zCUID1vpNMPfF1BpL1lIIA8m1nc8B2JlPyTu0KOqCO6
mVhailvtU4ffCF5VqVJHpalIMhXPdxBkdORCLX1upuSwJOkdfDbD712NzILm1XeAC2tBSpfluC33
ip0UalYegVpFvUbF4jpI6DMHM2RMpF/XkB82Dpxy09H/D2x2zkSclBAAJDhm3lXOfE5Yf8wrOu2z
Eit5SKkKC1BSUTi1kDEy4OIPmo1tVaIknST6yPMTvnyZLfwCOE5pewcRvZhT40co9rgP67yKCe3a
5pgupMJd1n5aiseMy9M507r6x5kJu56GufTijq/WK/Yiizbnqn+60lDutc2nnNDIeFMISk4AEdIq
0sj1mXHz8Og15L2OHkp6EPngTX6IrrjfBSaVWirQxeYAHgfWCspfSuAuKOlljjWH6AAqyDi63r4l
I2CzswlnBFKrP6cK1AZ/iPPhSJdus3NguQ0WgC+WZvCkk1cSYrUNXIJmGs8PpTrWSHm85YlV6HIN
5Tg7osWl9WUuSeLXEKpwA65Wxjkr8Ko9//QFWGoDmDHX9YMeLlivNyHCaSG1r90QcOf2PcF31w9f
ulpQ944bMNiH0QmySHDDqHUpMYimCQ8fxLdflSHUJ2UmLhx8qlfFRGVqyLyddWh7ijzIVfTaIDY9
Bjijh4PVZhmxYrHTiic+kcKRxfcPCYycnVzXttWig+fb1deqg3LBX8XOWtmx0Fb8T5zWyO+BPv2G
7oJpKriDgajTbWM69flNkQLyxsFpi8/KGsSYB1pjWdF5CfUfXmK561bbi8VL2F3MsGCobTg6UF9k
dFy9p+7QpeS5KmWhtS91InhDY+hgo/WvK/j5i7l0FbDr9tMDS73Nt0zGK1a29efv411eIS5498Ge
hjflKi8/eNHNTHd64ZhAGxXg8j4UcXmlo+G9qd8gyjAAzJb8w/n2afte1h4WVx7lm8v9ukO4X5/F
hhmjpPAmmTi8j1EICcjh8XpKI3WY3Fp/NAMsL59chUcS+tcUx5rMHCq9bd4NIIS4HFrfTkpKAzie
wnjDTe1Nn2oOWbUCj7YW0PmKR/+BnmAZR1ywjCz6J1HtntQvkfgCcuortc7LE0yjzbGmp5Fw4BwI
2b45tg5HiEnNwzlS7fo0bX8sRTY8Mxp27DDPr77H8X8pq7krohCy3dZE1AF6rjRKO3i6ol26C+oE
3omuCvG8gFEBkCuV/TZgzjA+dPPj0UEqOp1rEal5J8eVUcS8NwbVAF7BtxiGjXrYFgazHmk2KEdG
XZV7Fb1niVQaiiFRYNfP1r8+U7DUNjLsykGjoghvPb4KTvFRt8R2gcPxvzS9YsoZU7fdCb9EoPDk
e6cCjuFUkX8FOpRC7qjLRX6QHNT+IHh3dx6YpeInwuvm/YFYK76MaNBXXuR4DHVVGXw1aWMbJ/bb
Nwlk85wSugzkkwaenZt5uwtYkuiKzeTPbaoKDYNzA4P3FXq7CNi6EVdm0rGvHNb6D2kGR+5002AX
0f0lgr/kIzdBy6Gbm3ijdAV6hKbrfxuCmEFFDRczS5lJWmcROm/PyJAgmkJDffb7TZTT1bY6yYl1
U5fmRaYkTThrkY6b/vnjMXkYgQX4KCVDCGFRZi2anhFl4yXltxKDFYDAWIfTEnQZM2jyEI25v0r/
uJkDwzKHo0mg2mgWtbLRRYtHNYrAG6NYr5lbsRrfnnat67q7qhyFWuKbqSETdFaQSZsBKJyxwQwr
Q/oTfkz3buLZvPCBnhH41xgW7l9BufPhlBbMQiJqFt8v9u0PDMAsBqOBHVoAblRPh2j4Q0elkbdd
5zqdEIgvnni4bwe1g96nU9LYSQAcMdKHzXc01x6jY91a4J2eYtpzdx11/EHwA9rZbcY4atuhZ9Hq
cp09waexS01sPBE0xM1jYaGvpcoZwWblmdVs9y1F7+8N+I5F+nrXfgx5f1tVy0w9bRPlmDenVsRD
vKBP3yNzcy/joQuCnc+/I/9tZpXkv1fGlGxqeSTfa5OsvK1pSTsAJnGJ4sXy7QoIZpVI9HG6Ji1o
BAaKFD+5nIzVT7yirn/PvO+JpqlfryKb0CODPHpMJBTVaAXbjdW6NRlonz7iRuXVrqryHHKNn3wX
aABa8Kgrj1eIaFjXQG47tal709Iwlhz2oZTJ9cpxz02OXBCostoxwm1tvzXfUrENUIhCe38+fnW3
jL4WSuc1y8nDuxxED7Zn/ceK5wnaaCCqzhykf1vkqhKPrxY/eHB6isiJfxm2sKWsg2kf+v9uAkMN
6R+L4hWuC2SrYGJAtBOQeln+nkAHq1nut6RdABRU5rqAi9uDjXE+g7v1QLsG9gIb11he3+DzuszQ
yHwnmbAS9pSKBrqRN0Xwp+P/GToGK8T1bMzkrzMMj1mKFwzjeVmkwAST0GBI78wstAt2LWMri0Mb
jaSaNjqXmmORBaKlx0vwNFSCo22+8XpV/6lq1LkTSqSlkWUihVOcmlYrNTLrJzNf1DCFSA8+iySt
GX4/I2Q2uXDllym+9h+qZv41puxhKk1hmlqks+JVsTbHe95q4Rcw04DzAz98S/tQCstQi4zWbkcp
j3gQ9Bx+tcq8LAqK1LOdKEgXl8VTsFefcFXf1W+5BV+qd/Z0fLsSsdq0FclwuDHK5j0t7hqOQAJ7
AfLmXW8tJPr2zgDIIdVfXw5XYmNK54XTPF+g3zbMVog1DcBnN9prJreTZ1i/5y793X8bojJaR+mV
0ybEL4t3n5xJav1J8o3b+ORUFtjpJPMO+zWR/J8QzQ9j3dUpoqyntVwjggMgcliKkZvwlHhGTe4M
zN0IMgeIFu3ycvqyPFLxCQ822WOf2qj2w/HNKaHT6jSnmQugyzvKl3TvQpj5Gl4WkUudf6tLn0zp
gQyFsRAuWqqCnY6KhE6LGAn6vNfVm2VVwzCzDoSIxKicjCOWnOojjKIqM+C5Qqb6low8U8sDM+Pw
hkEyu6Ol3v3bL6oXWABB6I9c8+zxHcrjktTYWLmvXW/0+eDimeoGAFpG07WDCxARnwOJHqUeh2ZX
45DN/NrT/I+aryhOTuwWTa4X+ohcgscDzSa3Wm4NxVdGO818FRbXXu4/9RcwGXqGS014nRujDXSh
IJXJFIqaV8XxbsrO2KaLzUqjViqnPcC00SRd1DjzbQGMi78GLz4nNzQsUl0sU7t7rZquIl5h9qOn
6sCBkPZWrdYsJ7vNCwcbrCfDfkgE5/ADKIhE3YUP6IKCiucCCpqO8GkcY9YezFg4p+Fh1hXb6M8C
lkMCw5ZHpJFbyDJtd/oVw4/f2Ysr+nUSj1i4EMjGnVwVgHUkYbXvrhm9Hop9ii6BLDIi1fM54ZyV
89l4flkvXtOvNbLFU4ClSIXescgHdoIR1SF8u0jDV6cv5V40KvmpebUukx4EYaRbMyEqwcPDkpeC
rvclsgRsuqIwYjLBeHrorAEPJX8vKQsMuISgVuteq6TP/u6Y9GNr0Scol+1A2Z0+4+57Wks89xkR
pJ1rXpqtyOTwmSDJi7Hqfk/sFR0w/mUwEs1ZSIiAWqPnkrharpMRIF3mcwpCcME2U0v6gQm3GlwW
QAenGkh0tEhn9Vy3QSD1s+tfaN5dRa3ElDfgq9doo+ffCyCd/LqVC1zuOPn5E3ODWclQzuyuOT5b
QTQQeXOi3fArLcHMJwkotzMthJRVp7zCn4EVbPO+GvJQwYGSd4rOGeDh6HY1gR3dmZaFm2FaUiLs
R43e0FYc9rz3Yb3oU9U5z3BdALPdP+IlpdK0auZPY1zr4q4Bp2DpaH2OJpE0Z1rqX/oi0giPTvLD
Lrl8NPToYeK4RyMD8yxUnkdHhQsU/jfWnYo7s98v+zFycBkIkd0WXoreppw5FYF4dlWlTn3+K1iE
F1CDVi3OmBaiClWrP0Z/Z5lb3795juEP1GPJ2PG901ecGhGYjt/a2G3Ircn/zdczNujLK/w9+eoA
1a1LIomx6DUwtyVJtYgpST9tgjWzsh2Sbe2OPcMq8UkxllJ6419+Od+cyWZyZ8PqG7u4KB+9ckOK
JFvdSmM/Ie93QUuPGbsVgZkTCgU+dRc+tZw9N6sjNaBc0fFLcfUb6oWEJepcjjzqAj0a2M5TaJ19
dm3JHBptAmrEhpqAHatZeoFubDVGbjRjQWdN3K5CfdHIwYvcVxVCa5+tV6u7LudsSoDudVTxjrOJ
laEeaA2wRPwCmBoN4YPpDdtYw8Vp7eibsvheGRixHlGkrOkHwhz3rc39ea0d33AqlVlh+ZKCzchE
Nl45b6zEVDrrZONcT0X7EZ2AS4//GwdCcI0vvNCQmjTOyk8wUEO440GX6NKxP8c0kMYOG2W/Oe6F
nINf4s03nuv/HxXQ3M7l3TZcIe25P3xko3q+sT1mx/YVnyyGhVMk13rPSWOCNSEBgTUiZPHEsUn4
khOzM/yBqdt+MyAskCOXVqtapwUgb56XVey52Mx7zIaM2J7WUPycymiZiakmTCgyaa4OntKqpLYS
4Z92pwi8034Mu/chMIT0wKEf23IH9y7hKBxP0fpgg0slj8a3HlqsuVXONO9/LXvED43YMpKN1Hy7
lBvejTKIL1XNgasQ4EMTIxiu5Bjp9BaaYBEFQhLAgWmVGgGIygs0Yu5x5IoUSM8gbPgXUVGVqwPF
jHRjuQAtzFuEnyBroZb5f8k4cov4kldQUNG24kUyheW949555eMWhSy/bTQMgRPd6c+KfitnUM0R
52y4viAFeXQYNxwAy8xNNH7UxLQfRSOUI3xBe/HKKB5npvImOlJBYL646woPRBrk/dLGgUDkYWH4
pxt8fNyn34LpxbYsPJLK/IDtHB37OlbmqA8aAhU+ToSx6pA5k8GciRuWbtlS8PQ4qh/SOx6ogIOp
TwbXMkDled5huI9i1ybZOx6EkfMKR2oz8ns5yqf279gfsXmN9iSFNU+RFMYjnhxxbP14cIn8VszB
Jz0TDla44oCuTJJ7VlzL49cRrFbPANPk56jOekPFOPeG2ooSdV42xgEZyLb0URKz+uRGE9StkT5X
p+/AWV5v7R7USpuioJ9FZhnIOyuMR8MHDqKkW8A8rtkIjoK7Yf/f+cFwXZlg1xz/ntrOg0v5ETLw
m5VALvssFytFHYe8kXOZUSipp6Lgq4Yv+2ERyniAK871sql8r9JUFcXPVZcm9WdiYnIzU4Djh3GE
8rPHbM43/xtESHBH/yR3tQUFuwMJ+NeT3DrRdiM+18B2c61hPJcaruU3GInMVz95sODN20aD6Ncj
RFpvfoF50+pYCtxvoLJrjvs4zCbxYucxUrptv3BljjeB79bWmR/bkorkttj/QB6h+ZLackFh42gW
xPRR+dHlUjFns5iBeN2rcZlzsnphT5yoLB6W+DQArnA7DpHJ3xK52A9d0C4nukrQt5AsNJGhXMfI
qe3oU0OFH4rmN8WZHVX3sfEB8v6qcxUdA0AVKctDCaMM1LsRFsFv7SOji68q59tuCSCjPCyyD8WT
Ah8TxjiTgcCdgQBwSuDJ4H3+nz/pXbncdAVMl8EeeuOa0+8/0liGhRA+ccVZxLPgkkkM/7xLdJq1
GiEq1GvHjJVm7Bn6AjqZp3hI9xby9r5h4E/XiV4AKzacpGrR3TIWIvJxSbfoUXWbFdBs5X7shyQZ
qXe3xaTKEyEuRjBwDcjx9sizz8xMfPGQ8G+y1zGaTwQC6anv7fO3CCLY3pSdiGZ80AX3VZXzwk2q
bsByqV4wTso0XMETwgq/oZIYRJajZlZQin0tYzwy7Z/9dJDrnHyhHzTiqg1ZBwyZm07LFtB+imLy
BZfPmJvfoJH6c8wG8Wd8PgmfSYnwiLoFVZZQl6Vi5+lHZnfaO1L5LR0u6PkiDPT5DZHsarwpNfhm
2kyhdwNfcZE+mzXrhAVbAHi08l6wuCZPy8FdoUSk8Pci0FyyYBq+YHM/d9B7aY/vnv2FN9l3XyZ+
+rhdwBmzO2HnGVCb8r6XhBTSX2BKU5zZPmiQZ5Er83hdEDuBy//14h5zdQlDOUrppZLS0t92GEDq
5B7rFwN9cvjNKhovsUo+TA63W8wxohBd5Zves+5PelMSxwPHcp3BCLJ8MhK/6vb2wv0pPl6BV9DO
YpMdZTiyZ/+injgZd86+/CjcQHbrnljCroddG0QfW39ZpFuVudsaEijgPIPqyFg9FZ6jkkgqYaec
DtJ0Qj8oilhYQ0OkiBBcFy7z3gRV9Y5hjkmZT3mACJxlRCEVY3ThzXBomFyiD+MTTstvrJGp2VZO
xXYIBHHuQhEk5mAYfhDsN5+2mkIq5hXbBhHCa8oA6p4CeK0twXq1JbEWa0kzix2hj507pj6DYdIz
WcAmyYJhcgqjVmDslCgi/hjetfwwu6wrUi18ZknUG2Dm+VgCvs15YxJZGrNfYmkYnVg6h7/VPqW2
W/nCSgHbBXtGRppoxqAj1F+eiqgj/sjWBULHngl2aP/p6e3RoeTIMpmOTxaNMfyWDCayeosdv3WF
kfCKJg6rGyJVAxX700Q/4vCTvDMvxh60/7ofwZ0GKIpeFDsOJGCTTj4U9MJ1gJ9O4ZcJDh8C8lES
7HaemAWcx6VgdtWVQ7Hin9arBx9bp6FkxQG31Gx/G9CDBGMVQj0o0xXpVgdhUMp+n29WPtpuLnGh
dMvFqA9VWs5LT0dCYGsgL2pZOjADVeqUT3WmJApYOLehd3zn/rPUJm1fx3RFiLNZjEog7IwpX8ZC
m1jQlqFnGWj3LDwhi46nV/9cZToihgjtx4EA8FaZYc3oS45K/PvVcRDYAhWphtqHy3zbAppIpPYK
8go/0OdMOOYJepq0HxwPaTL++00RZ/0yNnzkMXmDgGgOZ4TVZw9Y7M8APpHCTJDK7etW1UiPF3yQ
eMNRE+oW3EUMNEgiVsipwfB++APsdkbHWkzSL/AQXV59AedWFz1MXtaaTmVTpkoTd1JqaN/t+Z8a
R1100VIB4wqQupiuLbs0NmzesfmJbQarfhau0qdAWXudH2CXj2vy4ZW/wuOVbN4RXYFsNuQTFDck
Cedrym2FihRWPcczxF2+BzDuCFppHPkRFfVttgbGCeB9EGwtP9RUCR+crEFhSma0pFtKqNqmGFNu
F5yeJMqHrTJQU2EpH9O8r/RjqXm9beqK/4yblVtrzCBDDM35axPPqpt8Z0+aqfzzbGiBrLy2MCfE
SOx5vhEqncp8ulVk5cs5IAfWxGzn4tYI8j6peus/t5pMmX1suzCxg/ciqdZ8NOta+Ss0rdQ73tKU
ebuOBwVZZz92z6YLczXH7y1NGGaLV4PHmFOwc73XV3uK4P8xaOGtKLrkYyhDooirvATAzqhcrEql
riJvnln9EzzyoiZ5jIDTBLVH9RPkMA8iOptSlEAykM/srFO60pitc4fzSUQu16IsLyVdAXXugAwh
8xkF8/8qqW55ru5mHLOcpay+I9hojijxnsvTCP5kqeChyCAG52NQEYyGS0snz7DIRg15XBROWR0h
sVcWCI9FlVcRRsaaVV13AtfLkcnvgkah57LEOvcwSHKR5tWbO8ZRi3UGnF/r1e5W65oJ1n/JIHLW
qBGzIBEjHbay95bW+87YFwAlFuUWUlXHYibbvwZPUB+bBDDX4pvKU4fbXPAbfch5xgAd+yT4Wj7L
0cyai+aS6MfvWpoBc+VPz7ZuZdC/V5aEx/sHyZS4iT7n482CXSD/cbLcHFeSqgL34sRtY+5/EmWK
jzlGUNjoWAl5vkZczvWkTGpncNJOjVKieo1DJ9iAKDop05ZioQZe6d6xGfl4Ms73iJNVJ+QYHcqo
B/9v1rruyiQaZrbwH12IjSQLsCJAJa+p3AuNUavHA1NBXOqdDnsMYu06+zjzQX32ggAHCfbXJ31q
MPytq0KFV8/RXs4PsCAk87u74mHji61cucPGHx4aXRuPPnrPeq70R5dtdh6iDeIX+A/AlMy7b68W
WG2nWNXtH6NeLw5oy+pHYMacYbOXEsEqJyV6q29kMy9VuJffobDH3858Tqd6lExJ9zomZCBXPIQy
zUAi2Go+hBUXYDVYX/+LEWw+qyC2v108jHCkMrfUXkWh6mDK5v7hivUnTW228IrBn7v+fiGKys2A
S1a90DJM1HpLL09IMiJ8V633N4RqQIoZ4mAhWvHjrH+ZOGBzMwYbRJegSZi2PSiRn3Vng+tWo/po
lhojwyVKbab180wr03CCQwk2zF0WMVK3BxQd4tmRyhHDvaM+8Sp4tQed2tHjL5YfFvgNgpPLEuKs
IH1xJsP53zyyzZs41Qub7JtXBwen62+EvnldmWAAumuSdDhOobI2k5Hts1sVX+RvigxZE5Y/Wrd6
DAevmKv2+dZjEI1wPv86nDS17E93vymUcB8H5tECK8Ljhrj8tyV2VZhmhh7N/g6GtwU/FhgyOE7B
HxC38sKl9XYrPTesXfJmH6rECOFINmjBo92F2cvQdG1PMXfmptN/9nXyYbXNTOaczjcnyQWTfCJw
lA7t2xTOISIchbzxwCmWmmsLsfOjEBea++2+7TpmJ0CD0QFrXxgZi4cCNPAv6+JwdmSHGOSe3FtI
wZTEIvYOgiEr/0eraORUNVsydF2BxdT/hqDgnfETzzjQl7f6Io4oXlDma5s/RmUbHXyJfgikYIDL
/GQaaISU3BEeKKLyzEUbmpm3OOY3cBp8Dtw0up31FwdNvLKbwcm4Voo66pKPYmzn6bUbi5L5y2nc
GIn73LBe7+Mi5rxb6ZNwsIz+EWCD60/EFvL6UfCXvo65nSq774oUY/83h1YX82MgNSWywmoCUKFW
P81Y8FqmX5Ivbc1yihdXT58voT4NJWXAHWomR3b8D/02U1WgIgDrmawU2bjDGGO6X6jBSPn/WP9P
th15T6et24wWExOuHzOlGWP0NU3hiotQ0lLEq/mHBY2kk10vuQOJFSGVpuUqswH+Ql389H5EGLof
erZbwH2JY+SYO2F7F44KNm8Jk37f2NF8a8v/bmf4UWRgWhZ6TcH5eMC/BdWzVriQzDElkO0Wma6Q
9ZKkJPtD51SU6f1xqNTmvIwtIkbDcpGqLHiEk3uqEk5f5ws5saGW1quYWh674cdQL08QG0C5eGmb
96f7XBY2oemoangdXwSlmDK7qZ9IgLOsgN2xxehDeruSDgaes0JuyJ0x/0InLgqCaLig9ZnkxJkh
gBjGH/TY3ZjqXMDr0hjSb35XJwVSQGCqiDQgNFc3praxFeyg9X8sFIDojly+0nQp9Qf/b+2B/kQF
IRrBtjbo/NqRZ+CJ1DJ7JJbsxuqUt8g/V1huRk2CzVI6qK4GsARyg3XXePcosPRZjL1H9KQTdvXc
q8j9Xqv4UvVZ+FOdRHm6k5YFY5+B4fgDgwcQrejLgEkw1QVnu/1AeoicCZWBvSPxXSiijhHTwzTT
XDb+TojxqE4LT9mm3/xnjVebYZP3H9qjA4Iv0rCPLQhFXiWFn7P2DIGsfa/ROJ/U8cnYaX0hYTDU
u7nOSL3kSHIbcZ1Mm1mDHZMPRGPJ/ZewywijYg/QtOW+5hhw1ygvWNhomM1+R/FgWFK7ANqrOUr/
M2JG9xg4ZugbRGhpXi/45ED/tsmG+uvW7alJ+wkcM/tzAUS6CZBGdziJUGwUbjVueCc5a3xDwLWh
chXaGPTCQVQEWBWlulS/XxubfYEPUHjbd3NWcQoPKERyenS5oqIzG9GuUegrKSkOeOKZJWjA+qQK
F6dl2dwGiZAugZeHEI5ReJkK/OvSY+lUg7bxy7K9Uu6atnKZH8JVAmTdJRwik02eT/4uQe6DJ9IT
TMJT/XzCxtUjO4hnD720vUp1EUuHwjjKIQ1NwGTYIEw+dJv7lDAJZuKCfy8GzzTWxs+HGFIwCiZ2
+EUOW3oYqgTuOcEqJ/YV2g1yEiO5gPbMDDryHTmffrAy2pfxqdU4dG3+jmpO2/5NuDRwuqtUZNlL
FXbTnyAeGO1J998AdUoMPs9x/6y6zPzgqZ37A7q0JkTtEcDVQAZQzEgSePmD1drGuDVmhNVm4out
411KR4ffXsWX1t09phuHvZqWGJdCzo09dmzkB+dvKX27CjIViOZgwky/M0uxISnYjMKZ/MCMh+DW
gxcMhoWmFFYs8vRpdNFbO3dKVsQXa2lU10LpysOUBEmH5wbQbQwssmyKQgBMDLPWrxohaeWrIXJj
OBPWQybPuZsPudhDs6xUIdfS40kxCFtj7naAMCxn+7xG4lMSNJipPJ5xkElt2MXj0Op+MvyRBi0O
y6H0bBOZOvHTwqpnr7q3e/uT3VVqUWK6WNOWZxRGQCXG4SW1q52d1L07dJPeTvHJR2sWgtmYd7D9
FJYjRIJxPcEXHGgYs3G5BS2XyQd6MzNDv6xG0QyLcQoeGZZUPMLOpBPybZ8b1kdNIrEX7mb0uF9Q
HVFi4rh9zX3U0TjrYjM38PITROzX8QcjglUK7VsIEaolVfipis57cK5BTEqyW6650KUMzadZb57N
FkBIUlus9YpNAInCbmCvxRIOGDFk3fZQItCVokNry6qmH9kLo7M0Zr7K3RwmQe/srh9slvbnU1C/
jFdw0ZMb2ErOWhvpYZJk1w6LLYhvfR1EHBDauK2R/lqh9M5Epy6I70vjxT+0gOClOqmmXKtOytog
mNXnrbQMGBAJPAI2W1jOP8dII9Sz+JPwJiAQwJSe5AHFPlYb7KdKrRfTwTRk2vAuBxggDvAWVZhW
rvvMcxtBhquuv/wsyz5r5YgatcAt3sFn2uDzyJ1Pq9WLuPIT5CdNxHicjZLE731+qm9ww2S2SHi3
lkxM1rfvXLXPdCTngBb5k4MrXqwc85/UI1speWhvC6kkMRyyLtnPB+/p0P/w9QlnAdWg7InWb4L2
BglqmZhZ5GnzxJWh7PXBACTox3PTuYPAd4Nk9bktUHDVlyxQeF8JXzcJSeMVe08N75lTlTqC/h3F
e7PTv+0Px2td6sYNCI7/Svt6JWZVyxDL6Tpe35Psc3YHQ3wX9HMQCbSvoHEI09mMHx+U4vHrYnER
H6qGA7z/mfZKQg1KVzgJ3kbVDs7s6YIyGb75gBQ0NWfyoa1wyAJU7NmlwkIuEDpKUcaygnAo5s48
WlEbE09RTVvfxFoNr61XIrxz8iaVnkPKskfKBZ7D8V3DV/Vad/dshi9YtlEGig1Ld3C0IsuWeDOC
W9qMWDYE013cFoqRnv/IAtA5pDrCidJEe9+LXO/tGOBJXd93jNSSjV/Uy1oSaYb46xQincD+Y7GT
53czug58Bk+bfETSZREx7OTUEPai7EQPiDzEZNMlPeXF3BsCWOY8W0aHIo9ButNG8DvrUXhMjiRn
M4CEe+z4nVG21e/U+G1pne9iJ5/1IabUUGHY7dxip0QgBDqwuQR2aygePXBM7crWL2WjH/oYF3sb
ZcrUrUIy9+3wibz5nPvmW0XXQ2UiBtrdNDsMDyGKB5fIWX3hGsjdA8HBE1k4vWod6oZJFsXgt6Pc
aDE7ZOf6k8FlEa/EBQWF8M6RZMBbQf25+E0vDLp1wvl0EoAtEkKiqNNWLEEPeXKfSTi11/N/oxQ+
mGXawTKdnWF6XZllEiExdh6z/vyIOSWgrOFya/jBmP6MqkjWKwKtwzuRU8sqlomy3N7AJwLXg7Nn
5DRDCJDCXA1QHKBh/e+dafWgNvsRAFDrEPPw3SriA5USnleOlZ3j7DoKx7H/XqmLxheZ5CxSF2AG
SVKpGVhSRXdTIlXuY9N5nvGki95dYbdqj9/vZIEPZGhfUaRdHGD3r70C/cqZ+0RvUxsn6CCcdizO
yoannLAVXTZPjwDPLdZxhr/npMcWeO2iisKHpR3kyZD7evUcaYCIHuVt1fwdiMlYh7EoZNiUMSPQ
Kik1OIRDZpzeRZaPRX3CzeoqyQiUgp2C8j8PukKpxusU0b7/UV014r3OopOBZSldNLPHO7hlGlow
ezFQr389xNdAmVEjLRB/A69n8uvxmlrjurq6xv62aC+PU+/DUao1REmeU7werLZUHNIwYrrrJYcH
jGEYYzFtlV71Ur/9G9zmmQ3+SjxhsnRfDxAQYmJdLWRZN1ZoWEoJVXxUi/jPb8UEgDa1xYt/vM2O
coLk9h32geyciQYnOkWVSvZJwyeZ7VgjS+BRd7JUbnKVIAk9JP9mS0hRCQVT+JHHtqtuFzaU4SWf
uV1fQJHxI13b7jRF0iDLtpwnX3aMwWhgFFw/PVKCduV0FpxY+8mGxymxhgtLUBfjnWG406Il+hHA
+nRUGBIYm8bhBemEZt8EfLE2v15P7JGKzcXkh4hssVhVzP7LiItewOPl+jjVRi6pwkhbwzkQtlx+
aNTA43yfYPM2N/uZZblcsrChIjB0mSxRF988j3YVVuBkmHfCMLifuhdN86hKVeHzbDa9XQk6sQ/e
TiOMLBc4dC35elSdF1JzJXCAjL4/0r9voOdwAp3y61ejg/+sy1oAjXR3QrJc2pSnk/jk768QIi0H
GEWTOcj37jBfKQflMevGLKJXLMAQdRGAO7UTIoVNihCoi6BZVl8X/nnTjnk45d2xCLY8QIe5bZry
6kPs+sxEwZ1CtLx3oxsqoCPtNz9gT4VhILQf5XGDaMALaNeWGYPhmnG5kToBGBIgwzTbEJgK9nEH
85jofu6VUyIG2kF7OiLvdC9LDKCcNg89R+gHDiK2pVm4pa5dwLn9iTj4cmUAA67ylkUl0i8MhY+e
88RBIbL8Orwug0mCftOoUePnkU2NM9plagBOboJJEBx0ZqwnXmmccjrvUS7g1Wdk5kNCAl9QI9jt
sZYY0xwFbHM8ET6RxEg3SdavNTkQ/00B+lHlojU67sZVnjw9nghd+DUDGPYiwjTgSnDvvN8sdgUU
dCCyDN4I0e3h4tJBpfr7Z1t4bp2ckcEmFpgQCLSrlAc11jmi7K3v+xX7uK3nBhZ4TkUQyKPZWf6o
dV1IEdExioEOqt8t+QFbN/HmL+Wwk4i7QwJ3ZhMfEOebo8VJzmFa+hOeWr0meI3xhA1VAEnmiodO
rhZQ0oiNOXJRaHhiLdB7KGsyCYJEoGljb6jRK8qk3p01LwO5odFpGNS7eNob66tfFR51H8fmyNHs
J/6tmA2xrWsRMxc070xYpz6XnxegOc57AIdwAQ/9qIGblRfxPli64J2tDIPfB2Z1zNBsgISKpWpH
6k4jbkCXnpuV+Hijihcmi7qUetUpPIlZZ3E5kzyW+viof8LpH1WVzwBzUDAnxa1AMztB1etWYGrz
2iDFA3mcd+cG8/Z3VvIVCfwr6GyHIkHdLN9PjtnKImSaXwdb+M0P9MstkA0qzzj6/Y01IX/nCIlH
kSrN2xASpAVPnlVvwRHvjXrZCh8np7tSK5I2+zKFAF6nHdbtwsAHAzHN6V7ZlEVt+mavTgQJWnc/
leNXunXPs485unLflewNmS8sw/9hVAwBjR/VoiHqR9HNvGxnUU6BECdOwfj1zBOOtBoEA/HgKOQG
QYc8Cw02o7DjS+kZsx0YK650PFpdXheeu8Cv/wMsrDM/U+wPEFpyMAjP6AOfBzhu6owkP/WXqra9
iTesNeJ4yP29TuMCEnCmcRbUEBzkfHUcarcgpqnfxnjxKmb45UvizmEreklxA6XbXLXThVd+BIxE
hofAdUtsDxC26y4ez7n/FLAcAhyWyskqAG3GH/ytKrRlAcd+Y4Wprb0wi5JNjcALWsPY9nsQABd+
7MYCYelu60yzUxrUuHI1PEgAjjcv+HLeUXcnpUP5Bxevh0b9yz+WmLQtW2p7wDroYpyby7chTIk7
lDKhFTO1i74+UGn24PE2Mumpr3ZKdAom3VL8JYel0MHNAtOjazqGBT1TWpPhdPAzH5b+pEVYga7w
N3++SZHTNcboHMogi2JtC2b6IdZBKE6iq0hyzRtjOH7RuFNL+YYXpuPNch+5sXcev7Kb5JY3LjSt
gtZJSPDr4eUM8GEu7uf0SE15SJeOB94tr4vmFVdji1sdsDyHJFDHSCfq0WyoN/bW89b4JdBr2RH4
Gj04iaIGtJtGLGFHPuD2CaMutAwXIf6cUsv4QREwOGjIhCV37ko0SVb9PQUwv4K3jB8vO3QQoSke
5I6brkJzexgJrpRzTGjASuwn3pRJPlY9FSDg/b7XYhdvfJQi8SKAp4pFhVy2zsSJP1YPJpiQc37V
XPc9LbpXCxRwCcjWtn5/vrpOPeud5KC5vIaJRBKuCTA9ZCYsKMabTRv0WtlQlFLQbfHlARevTrDQ
OHFqKCd2ZnViJiySSGiIxqskX3tyFUfc9mALGl9hmGN7njvneVfwtfQlQSR+wpEtmuyyyag0VUTt
HqLbUQDBRADgVTUjcuo8lw1U5ApkSfxSgECSODwEsSxgQVVirO0iXNm57JwZT58Y6vZrAEW78ReA
Q6cLttzy5JMPtjrUmb29HLKNVjRme+lWAVf39Atj2dXHvgI3ertL6m4Q9V8ulej7GuXmYn3+7Kxx
Pp4MOq+ofOJRfQXBYTiLma3Zvp7Oatu6F4GbUaW4cObFaJZS0gmbZL9XU+Qv10JWdjqetYeGEo4c
/furjVGnvvGFWeMovluJvAVgrjQX4CUSc1t7q719MkBNkKfh7WdMTG0FgD8ui8k968qf7spxfCEE
NpBC6uBiP7FOsvjpgkDLEga/s4Td/0Q1FMrDsyBp+GDrVON68fCH9IdqaJUDfzpxcGuWkTDjq+8r
DV+VZT1a2DpS1FsM560h/JO21AvuCy7lR6mya++bTp5H79UYYVlHNreb5mJoaSigdwCzxjR5o3zu
WWKa0z/OannxZ9Y7/AClk3iBRMDmAf6RuQ4jqac0mYuyi+ctYYPLNxEZe8wBw+6Xe5m07CL1aL0G
+VNYiLmkU9rtN1V9Ccf2h1yV98jMdNDm15kopXlRfxK2G9dueMiTb6kDTP9S3dxl9O4g5MYlNu79
myS465tbJVT5W89PzhIFGaEw4R6eCe9JQu8w6h/SzqudDiRXdtogK30D9T+JNgwY8B+b5oq3xCyg
69EbtrJc5s0oPR7T/VA6fmg3YJ7iEdlwpNoqSTliVR7iaEeyExo9NO10bCXzYqeCjTcQ9fAn9Nbd
S45U9RpCb2fpt0cHAyUyNIeA6VAuSrvd4Gb/G8ZrMG7IQWjk/X/wz3wPW2caSsUChGZcPReBJz9u
T9OpeyXNEC/zipIS3EGhMh8VU98yrMoEmGsScDPNklrVZj/w1pPV8oMmrbCNNa+ZZFS6KMtpj/q4
oIxm3FrBGPdaH3agJHMYAmSRmlF09chygf80mu348Pp6vXWpMPP+WFXc7oA15sSwr8hBXV0Q0mLC
pMQbkDPvQWZFw/u97ihbTt0rHGeZ5yo8rH6HhxhnwJy/4IzASBenjW1g0p7hZQfroRxdATUKuMPg
vjCvOjJYJVLxmHXZNFLw4qXMUNY0/UymfZJG3RQbt9YQMcC3vfMDgNyk95X+vZp7gqdBFqBv2Nl3
EdBy2Oaeb4BdKRdruWzg90DSvzXcIeGe+xQj7a1zItkDkM/HLnJpWOCEcmUPkO/nr4O55slLW9R5
K5jBQGPG5BHso62sxcAGjukvixgS/eolDNYYnCes8L0fjc1qS/jROKIwI6CtwaWXGdZZsEutqXIy
BhLk2yZkBemMZh89AFxvi9WZ8tbNQlwlJJz5hdVRhfycPQC3W87Ye9RN3L564mEpvaoxk5/UmlBK
zKKe5S0Yd2ZEJ468aRSySPpEPdRHkMzIYXO7aQNkIwBfuQJjfFvyFlaQJxD6MsxkQG4kS6TaCxev
hrLsCMKGar57urM4yIFP/6LsWwFno+18Etkk0OAUExMDgC77qqHWaSVwQHWcPvBFXoJ+YwzfG33e
1AfNIDARH/95lPZ8nzOJYY9ezr3brk0PCnSK8Qs/sAPDsTT33IAst4VBTY4MdBhEhhDV9y1qnVt/
zew6OrZE2enD6cRFPaqCvSL+iP63NBFG+0sFMc3iXfp56OlAKlf8Jso2A0qkeRrUHPaC7Ks8dUx2
QPHqmefqiutqgJgjU+gXEOHLSHKH03VeGi2hU9K2ua/eFTR90M/8LOPnMVu8+i1wz1hpvUCpzupK
kLsfa6BBMcuGF2kMBYW5YNBPF39dbLZ7d52gKlPr/PSKycLYWqJ8FVkILdjb6nvdEbeF4du6RLO7
WeenEIkL7tObNjVrzmvjxaz5SYJwqIh80UK7exXEC1dChgNUoCZF5Q4pxHv8thkWoRawfSg+kboo
8IzDF6Mlvh8/TPjST9tggdGKqlyYMaLFjPq5UXwTZ1Eyw1w0G9eu/rBfpw5DoNjdk5+N03QFDWSG
7/EyWmjunshUVpcJoSlSsMD/VZ8Q3hxsG+ioA5G4cMEIX81hQIPugs8olKq7e3nRHt6g/znKZNnI
u1Stm/sofsmgzD1MBwjAunynBFcGXVpQ4fg/MTA5D7bRXVmZqRB7aAeKVv5MPMFt+PPRzJn2vWCE
maGujbMySkzsGyDupcHynLyoMicVbChQJpuQnLf+3xgfxgfDu3CRg6vPLwyF2aLppQ2dtT59ea9V
euXcJuQtPKagKScWY1znTOk2ABQd0ck+vHB3bTvpXQE7D/CpBqyhz5KIDOcnEDZ9xzJhjK8CldVx
phJm/QEN5TNzGTPPijz5JdUSCkABXYtjvwmcLzz/qpKEoAmyi2KvCRLAf5eKSp7gdJS6d/4XL92N
OKxqPFMdR0QGG9G92CUSZVaRmyYam+8jZQ3l56g3MXB3DmkSAclORSq4kOmeMx02n6Fh/5/xXlbe
Nj8EISCsxL3eeitWWkagTfgr3XYjiEB+P89l8xIJzmMzBTkyLt4RjsQeQLm47UeA2J9zGc1wjmWo
aLNW45fiOnPlv4MfatruGHp1ERTwhEBtgcMFdBMP6Ezb+gtGF5NOaoO3i2SfmQv+xw9hu/+I2hFc
GS0hC6Abov1PTOIsCdckWL/71YKMqbA2RCySsDYW6HZh0x6MqnO8rlmJ+M+UY5dQF1A24rq2X9n0
U7kk8qvyrpg6T606kniqKIvl2LHdfv4ocmRiIL34mxDftfsG0xg0Eav2Lc+9IhrN/720F7gj6p42
9tBJT2gPsS71CzzB22h5BejMDq3SxPR9ISKMcoTrB1IPsjnb6iGnB5CJWn6v4s9l8k22uepSrk4U
ArnhhqO33XILFkh/Rigrfo6PkRgyiRMXw+e/TGE5qYrO6qau/xVA08ORMMqGVaKpYF/e09o5xuYS
hpu3PW6xzJq8qek9jyZbWWbipiUzDGH6QNuw2TSWBQgsEarNgnlBqQ5e6TlL+xTcB9dwOJW8Mm61
FYIC4YnG500T5RVqDteN7j6K05JRHE9sXcLZhKcAbFaiU3BFNYv41gB+ew0z241UoyG5Dc12/ouW
EhsVfIevS4iNmRqO0fgRCNqCKQu66kv+CkwLixMrZNfk7ePY29QtG5Kx5ArsNXB6j4shN/e+lIwA
Ms3VsYW6V4Qj4htGC0ML/SHsRLWUNcblvn38RT7NT0Nrtpvnm4mtuar/ovTbb73nbQ1qBVIcFpyM
KlK2um6sH4cGHceZ8RS0B163J5O41BHD1WyQ0ZaV1g6rX1AOQ/PAGLKMU0Lw30fhxR9bWzWNBskk
VabV/4m5YW9efv61eyZQpc8qYud6IZxAKH/Q7N0t0tkWTPayyxTuG5M1QMVUJO04jdVPmxdZMtKq
zxtCLYjLNIXPpvB1gCSi/aGdQfhmUAkuU7slfhhnAO4MToGguDsrCOSlnFrT5GB7ZqAXLA7Z9Lqh
YSzTQYtnZ+PZacDQb+dmV3qgMsgI9W8FEwCRBbUyM1N+nfM7Z4MqC+15s/IWd3eBjxQAVi4XQt27
Acuw41YmHi2fQKTbbqRBXmM+znx8plq9m3cA6brUPUpM86pEoZhfrHMUe4PA+1eBqHslQZyKzVCQ
qqoXpmERpCDw0MXv9stvhDEDDODrCpWYYwkng2YF5YcW+i3lsvDWXBzQ1eUcbUGqm2LkmI8snUpQ
6XWZ7+94W49dECUNioaBWuQDv0vpojhaxrHF1+Qtfr4nwFlKT6FYjkWYl4GSW3g2Qp55F/1TVF59
rpaZqIJ5HKe1igkftgzOS7vehBcoy9NxugBug/BmbnYm4tKDmGpNQlT0e2TWYuHhPK3oOxujsydW
1gb6sJVFDf1rq2taNz4c7cJbxG1qvovuv+ho2Sc1X7WN45DjKwbz5u8OPQNzmSOOO5X1Q5E2W8Ce
k1FeLIicEjbmlHk8LA0E867Ix+QmHmkWIhPk6NH3CefLo9lzeiKO0diLgsYeSz3OpIgbiFovRIVS
cW1p5VaWHQYVlES9iFSrSzvvZReODyvavLgHXScsPIYon3CpWBwr9FMlp9styqBNTMuR2Kq05fRi
thtzVYlksj38k/CMSM/9rY4vEJ3b3exUxbyEzDIvO/B8O+ymqr47NRfETHwU1x1NdAPLfL1pb+wL
mB4O+t5DBEi90LO8+WYGrNxLCOLMhCRgSGCCvlIvcuLZygtDQUH4T0C4AzG5YNl5Z4/RvlpudZk0
A1mI0X4DRVGTvRDCHquH/EpCdhLtDT59NqisC4HgMR+fcyKxMsd1K2QMOiYmB1fEoEdKTI0Zd7dw
Dd0zqxYmLXStu/nKTKvQN0CIqv+/1rNfVxXI++rHZzfO48C081ZWHoVW9ACT8aP3oi4o0VWbnVdU
dYbJlEDR6vNIOHamGi5gGT4igMI58fxwiruwDzfllQPuc9CXprColuBxMMNnyXo+boxIOHvGcvgT
haAYn6rLQeeN7khqpSbz8YE1qriQMEueeWM4KPVpBFf+mI7jvOVDqLMc0UQgeKQgdZPnioE4CR75
mBRglm5JPcMVMh7jKsSJJ6fmguNd1b6LS8QzCdGIdgSJdSwOeQnFYnVn7bhe/LyeFxSST+8i19pM
cvI29Hqk2CJPRXSfi70tQdN6gzVnc2UR59sX7cXKgA1sA7dqP+LsiwHreQeoo8k5hdRLV+3XQ3UO
QC7PBwqh9V0kLJtnRAwxoekBez0e6zbmWn0wxf9WWXD861wRA5WhBZToyL+d5lGS8VhIw+9wikfB
zDjL72OSnPTq45tDwFXFMxYU511fi3AH+YA5WCpPujobBHizIGSTQ/DcSBZ9Ma1jTBUOtf12zP8u
KbR8alKMUEsh5Mf+giLw8roQncFJ4a5VsCn03Hmt3JzB0ws6DaGCmAWfeJ8YP15RzWKwQJNbvMtV
Io+sxsKaeoj+v5CCCf0DYgZFcyABGsmAuPkOzIyI1768IJ41UBIwaRfwU5p7nOSM4+YQBntuNUTZ
SUpC5icozax+CmWxqi6cxhAMZR7pw0tbzSbN+/HtIWWCywEfzh+IKBpvTi3mG1oIN412xCwy7vW3
0mB2HctLgjCSJW4svciE1PY/ppsY814mpxuzfc3zBDN8+FQoAZqvLaykF1Cfy+fzVWy+ui7qVUlX
LGhlRhhnCD5/KD9OjDAtgXHYvCeohKyIDb/RQqzdCeCv+NiPO4/ZO52kSvOmf/BJQizW0jWzlSCh
hhLAZk3BgWJrEjbIUv8qKwTJGjEhqEsL8AkwiB5HDphR15Vbhf3eSxK4VYAYlXRm0/MokUCdKeN6
0IL3dlLiFVDUW9biQJtDlJ5muxEmhc/lUZ/jr9cPxnW44SwVaHUgmlNMXKUI5wVUfWEnqh9vsoHT
fFcl2y6fUMYkuBOMI5A3qORnwMPFNiYDHBd+agBTaXAGessIPsyl17wzLXF/adKMqP9swadKp+iU
ukvXh6mlJZ1E3eIbSKOMHvSpSPZLiqRBuE6qNG4t+4AN/vD1TJNIqiiM2Z30XkhmEDKwXzVlNjDa
D/hzNSheQPA/7k9k7wqfokRQU/12QkCmABM6IVkV6qIvg+Ly+/czVIQh6ZukJ6WW+ict6Nms4NkX
BM4RTZDQs5fBcshrH4jUelfL82X0S5rwRYTIYNFRCM4Q0WMGEjNK1TxdwLV+fhhyRSu38c/A6aJq
gJjPMs7e8ITq4D+wk1YFk6WRDH24JqaevYzUc2A/fL7VKSMU6FuwTsC+uhPLkj1WURg9BnfmRfS7
YJdO4xFaDjJIh5u9fDrf4uKai6mqXx2/e3oAnwTEyQUp5qFoEVYMoPRLkCOZs40s4rx/HNYiwBrV
GTctNnFEtFQ3hMEGF7f6QU5kSkJ4n1Q+D1QV1WLTUkpDlZ5meQjnLCllMSJJIXzcNEBBwLKLwFpF
vgcGA1idmgPQHKyxC/J7YHHSkhE12MsUxlmOXKu+kkPfhcbyb7HaLymTpdHhUmDRYzDGKFSSRoUk
G+/sy414bGkvsxxIS0EhhflpnDj9FELI7+CjL9UKTZvgLWqf8hxwjCVm9CFCBeqBFBMH9MvcqA3c
lkCzKNDZNGDR8pY6G4jVAwNwaVfjRk2L/cp7ZJytEQhJGOUO+7h9zTzNbRtIXEPXNvhkItOS+2TL
W/C2Giqkk8ZOOMsTKxOnjiK9yfd+otHysvTI2+Ioswc8ywpqxw6qT3sBKQ1wK104jXDJTq7FVxje
+/7EmuBjqOSzRUVrAkkrRr9oGyovRm5v5LhDl7YGdiZEeYMD18rN8XwCvRdcM2Pvx3SKrt29a27h
GzjWdIx9/Him88UA8wkDdLjh2lxoWp6ImEetWgrHbgRxByvQlME4GbYlLwOXblHOwrViPnI9ypyT
r7tWnK65mnkpFYnliB20fKjoGydJHxJCNB2OcDUuTHMV7wY0AtnXtHEC84ceTgNuzpf9XNpiOgGD
VC98pXXgnuQF8A4AYn9qw8EIvIM5FpSXIQio5PnARtkY4zv5wW53taxgP74375tVkk+lxULCs5Q4
5Kp8kuFAe8V/EQ7fLHuFR2ynbk8iYQbW7TIRCBehbErqJMjki3wzxrXfCDXOxemlFLTgNb2iYUQp
pNzKTvyDG/lm4xab8dp/Yt+yqSvE9x70khtUCs/C34QzztQ+gvC1Sz0HfPvQ5rHOobk5Mg4Brqfy
yOx286kIThqM9MbZII78+0BglNoUgVtFURep8i0bkGMpoR2N69WoqpeN9OowZNBkFng3RRY7EjZ3
6cziLkhXfoVvmgZc5QdyaEmH7GGA11rU+lS06fSQ5Xxn2HU2uK6Xe5uSqUnlnr0YM3D6YzOjj8wH
xIYkgaBjH9B4fkUhss2xEYjJl6Xg4FkGxEm7vZtRr+42QVAOigtqFbOuU9s0W2gEiA81zbiNIjHh
bHwr/LeFRLVymCvvoes1FSdXVUf4F0NxGKeJj8wBYA3DidOmcd7++yvdtW3i+wUysuvc6iFNv2gz
PqZbOFM/pfc9GbPNwQ/FV2gZ30OmOmaXFd7SS9X357ppsrFW6dcFMIjCubG0qjtzvqvYCvh3BWwQ
D9jWKzU7J5U1U7BSzEKfAfCnZYDJPodzPKB5PltxbQeZ7tHxWBnOuoQKsaHhjy65dM29FuHB4cgQ
WHPIduBzTzWjG0qfYy+ZFm8fGH64f1KM4WnYcGXPK7+BQqVWjYlNqC6LEmGVJ28n3XCsZmu3kMl0
Mmk/cyDq2kNO3uZq5p06rX47UIFWp4ju6wlPjZT+1nbNNpqzXquWB53lyGjnlOwe3mYe9jvZvxQv
f87aF9wUGCumPiY/SS1VUrAdsbrnIp813Mwn5pNokAHtlw/03qKJDipPGpVPgfCWvmSBvl91CPoW
GzaBlUxAReJPlkqghKR7haXjujIrMqjPQ6+tZu+uKt6CkFAZgIz4Q3urmEOJEDWmxJybn6Xc0SsM
+deHE2Dy1U5ElX3iAy9Qa9dbqRKf/6Evhu64c4pg+FqO32u50jMsAFyfe7/rW969AEFmF9lfOBk3
NQqXlBosrhiWVLQjCe6efbfkYU7PlBv+Z0YGHS+JZ/4uXQv4abHc2lKEXplz68jfm+2ndYsi97tP
wU1BSypkQx/5L08R6wSTIqoWtnMfE099uJK8YmyrchvvE1oM+NSyR+Hekhs1+GR6jiDKOKe8kN+g
0dgsb5ECM0ZRLJ3Z5d/Jew9zZ4y7yqmLmM/iWgkmTl1AYI+Bq24Hed24Co3+wNuP+aUI9A9C52gl
ru8v7gflEChOtWuNUndz427mjc/hw5iv+LG5AM4JKfwJ2JIjMctse0x/cOdjftn24rh/JIM7J5bO
sFrLvpSVqzyXYtdaG/T+RsAlm8nbrb7o/TqUTgePcb27WPrBE+c5HPNU2SxqLKu9aPnIixTWddtH
2xljtTiFgox3OmE6d/qKw3UvUUZAg3CsH/SoVKcugLTxQeMC5f7Ta4ohZFBeuMqs2U5SuEp/OMlw
pqHIRVFF8CtmesW5TPrCqA37L2Nx6EothqBRYui+/brp8iJHhvi74aMxXwz5YzESS5l4TrrX2UW7
j457H7wvB2lFVRYr2MntiSEzb7M4yb8xdi1+OpCrN9iC0Wip6NCEdwtq03AjEhPPLeLAw63s5fXt
PFwJS7HAJRSuZ7BOHc2bVyo7DJ7vyWVd8KeTNrsY2LcTW2+7sM/9xcj3O7RmkzAlvLqE3Rfe/kb1
i2XMuZDIe8d93sF71z5TvgPGmID+iIHZPF9cU1dcoxckuJk6I/8H7uF1Tspg5YhJ+2q/6XeBqltt
sMbqHXwJ7N83JAdIPPWXwAUz6X0iDCdgEd7en6hf6McIkyrFNhQ0+FIiPzaIuxTh1ZfkCSdaE6nc
yh6r88Zj4GegDeAVCN+szVu5hdDWOcNJSdWmjh6DR6AudigB8oRpIPX0iQy69p7T5/WtEXWmQ5nI
yW+bIefLZSbo4sTyzUL9Hi62bc5jwc/vwt3UKs70CoiaWKTaVCp5XkswlbLT1QgQ8Y0E73uQciPH
CeX4V59GLj7b9jAy9PAgZwK/G6GpYrmij5ZE+DXWEPkYjqKqm5xZLTgliton4NCDU7Zdyw4FFJTs
UlbImsPay8PAMTtFujCoJhmA1G74j36YFUp55KGWn7dA5V4Jn5hvVYcMu9AseJb+ofxZvWV53n8z
8DQ9678ii27SUo8oVHe0LlCwcMVFw5DDldvFaZwcTrFvhHxAkOWKYJUungMuND933vi/nd38TWQ6
AM0MwtrEUB72CVyhpWWASBDoX7aEoVcF+JSO/HRdztsaxN+3JMxJclSXFOcKN+m6+UvW9B5AUq6y
CyqfDDwGWMzh/KaAVI24UEYJizjN9CWXKvmIbudqHZEm63Y/jn97u3cZiwcK/EhgK2lK9rieUtYg
LQfeA73ihTd8CljuJFB7qdD75htQpqjnN2hkF+tQGE3yx5cGHAej4DVQgPql//Jg8Ygcdwycw9Hr
+8rWkH4btQe7FsQBY2WXAndbah8E5C8y2O5JV+thvUe+UByMJIKUqOC29maeHQn+Ed9atetWfVW/
xbIUZr4RRTt3DuJgSWD24XS94jz6dLT1LJuIzYM058L4V+70AFCaoxhrYgNgLxp1NAJCMiBbn2W/
ahCWWq5AYKUEGIthB+TDnHRixr72VsNt3JDEd0Nhxq95DZl+lWxa1rSqbiOImgaAWqWzhrLxgDLB
uBmau+IBCpWUN66Z2RXp8tn0P7svT9Yrb8BSjAmVYiphybiT2jjwWdG+leKlFIhVizVclvpIA/9q
S1VKFBbiVHhZM/YGFgfjSsv60JUykuyztVKX/+xiUyR3wGn5FgKojAjLHIiZW0Zv7gGRMkqTleUe
BDAIe/0viuQELAI+oLKmkB8MM8TezT4qmWeU718NtYshiy5c5QqBTtVOswtLJmCXHBPn7ehorHNe
Nu0Q8CxPr/aDtfK14sRBYTdizO7gSmZuHnXG6lLFd0nz5RlvFBi6HXd+lO4eaoGIzMFsI/m26zAy
LgCAoKJjJTWnqVD2npXskgAqBPtTJp3yYw6+YE5WnAcrkiNZ3vegIxhb0es8jo6hDQUP4PsOVXyF
eSg8WGvISrXxelrdK2X9EUlHeDVGF67/SEVcloA6faXzeUvPNRxWgAPf0APtjCVJPASld4zI6Jr2
GzRYhPt+ksrXUFBzZKOIqKji3JYirdNoRHoXK9Sfhq28m3gwJrJot2cnC/TsuXLpPzuwi6biyfFc
NuFCy+a6m2oAzcVOeZE5z+GPrqS4GwVT/BI4/k5rKL/snO2h+4g+wjOkKIpKZeVR6mXpuFs38+uM
TZA4hVr89ycME8jco5rlpcarS8H8736LwXeZAkNZm/MJ6+UulkRgqgffMUGF5vf99Ns4ShQ+T9xM
tkgrtDpZn2YwTP62EXfYkrILeJ9C3SrZSpu81zbIRkTLDSUo7l7rY/6BwHJEZb71MciAU6JaIQIE
Y3f2vZixoaR0KT4mjTon+dheI/FFYM6RIlWbXmNOifidZ2sDAD1dTT1uNY/6cEPVDGI3BI8FDW7y
hQnkJpAyKjLHVT9gu9Wmag4cqZY5W5TQpW7yAbPiWNNKwD70uBSK5cUWHGP3b1gygLkJvsactgue
3rx7cWwJndAc4K5EIFiyiEErBqJIijWtRdCyCIYmedxI1HMo4I7cw/jnRxpSYnpSuoiOd68Ir6gf
FW68eBujo+J+Zs34nRV1fcUtBz8J536MJ5ZzAzP8G7yM9PlpDSKqZprIVPtxvyK1u89i47jUo0DF
/OJCq3MC3y28y0rbZj317z9gXWvWMT+BAH53lDE8l/Va0FW2v7ryioMbxYgQoZ1Dz1Qry9R8zdwW
GqGHlE1A62+X5ETjBbOGoLz9bL7N9AdVvnDQQcHKqz2CAsHP52TrOQybumDmUX049/SJLHa/ZrNb
0F4NzjqYIJq6JaEn8woz4NP69Bki0TeHF+bjAEwijEO7eSrpxlUpaJLHK9Hp8Nuoi1An5HZ7zDOU
XjoO9LZ2kBclkXw9GFBlFFAQ6cR0K94W4lLY0p5s8HXRxoCW1BoM1xMuFcAA5JQAm8pp+2rg2WUR
Q4MpuDCpRPkNCTLQcUih7bEz5u0pM8CLpkiXH9w0equOTZ9iHPkMNbX5t/yMiyFnmEskwdsmuQiL
9vJV9mZg4M7HzxEJhPd50r0uTJQgY1AttcweBNlqAHZNYbQWP5jeGyf7lV2GzBjn7m0bW16jwEfd
8I+PbL1wm7uDCwHDevbyqaqsc92rpoeg8hzkKYBEHLEnzt+M7/bdHm9RnF8VKvE3HpjuehphoWlC
CRUe0/liAbBM4hj0bPideW4MIzahWxgrDvfjIdlBGDxBLWirzpvNJ3i8KBPTRa0QQDGgDsWeDUaJ
4g6oUcmzxAkm/WyIoRdLEb+Xdnp3MMXSzUUXDBvaSEp9ZrQH3ajGsWpoPaZR+N+cmo2sMvyZw4tp
d13sW/CNAArixrP+l0QAdoV+fi5hUXPrM3ag3utXHpheQ1qvMljJaJIU34ihJqgxCBJ+aIVyfQ1H
RRM6V6hRBcPpWHFf4rQPZcoab2WKdlLyLOwRSxm4zE5QEVJ5JneQHHmz0vqlvM5j26UVlvSIITmd
x1QIzehJaiKaPa49j0KY9mJ1sDaxcBIlFULucDUa7WaH+yhnlTjh/FP5iNgZlDgcg41X4IcBHWuF
chPq76SJZF1hgTpp8Z/n9n6LVCzQol4Jaweo2wjIxyulZqM0Fd+sBlS0nvUVT9Swy2yknmgHEdgZ
TIXHsY8cJjO+C1iOPxXpR/C4Q2wW7w+E9/IvAMnPzEC5HlupbMzGUm6KTRxgP5L9FMB/2KBGVb+A
AObJCLKbDnSU5WoP5kMOOQAAUiUYtFVsgVkU+EL+uwH7LXmVeX8UOAd4bReKQEVhWvNVg3J5rmNs
dEVqmUCaGjZSSharItOsg+AYrIJaf81unZKAtqwbKjeyk1X54HuIJbqgBExPnJCHdRu0oKXRNNL0
7evYEaefx7pi9g0tXXAD/4VMX+Hg4ypoMgiDluFwrUpZ89p1D6eU51NeSVrGxRdMN8VKRnFXaoIo
KLy4ikCJz5j3VkubboSjeMy7kfOtYSHJTFkCrnIvRBviA9glNU/2awKIUwdPRKLCN4qVjYpjkX6E
Z7N9JFSB8vwG2HjH7IAORvhpMdDQSRV4DGVgCn3EBy6uNIRzK8lhgHg6IfNmx1Pvm9M22xg7rTlf
k+nleTN/qZjCPx+W1UnkS6ZBNT00YhMuigxo07Kv9uAA1g+Mi2WdagCaaZR94j0hozNyfF32XAx0
AWE/TIFZUQtfwcbxXNslLmSuQWciSp6+BOwnYmTErR657owXGvhXmxrMuZus07ct8mJhwY1nCzfb
nfEkip942+db947D+RAz8D//+GTevHGSYS4IKllz2PzeDi8RjhdcjA/RH7hauYyBcL60IPPNs5SA
S/pYBQ0ldqmGzdWxlO5Pjil7mG9Yumf7aX6Tl82OnMR5m8l3Luuga6662FJbRz7iou/E+UJBp0UE
RBYGqhWrNEUV3I7taZ5N7qv43GQ/OOSWPWBskgtnNKJwDjWrpt1jlmRpy9cp9BaMdCARRISc+UnP
WqRVDrLszSHR2KrOABbH0oJk54GpHbXXbEUXNewfWoq2kGb8paSmLEpxVibkpCDlHNpDf3UbwEWa
umiW8Iq0qj0lbt93WEy/qiB03Lo5wF1q23lmJ6E3Rk5TDUb7zhdJuAVQE5kS6Ve3BHxcVtaZVApO
EVWSd3jgrHCcjtLz4g7QdF0a1Z+aqzz8Uk0O+mFGY4xDKViR/x5UULUHi7BpwSqOnSZl1UZSiCwv
LNB8fYQATsbqCp+88vlEkhENoUc0/8X89ONzhWZe5eZjwRuafDhTT3vWIm4lmFULIrOU0xA8r6m8
25mZv7dnMRxnw8wOFI03JsIWBXdwyYuVfnW4OmmCGP+r6RsZza2sNSBf98qZpUh6tpe4WFov5JU4
k1yadtfhXQC5VP0FJ4i3JbKEy2edmgEKq2gj1y2/Rhdv3PUMPwQZths6iUNVlElfJA3UQ4e3Dfdf
ZLWOfP2wY1U2/yFqSiP5C5ggj3Z8VsPsmirG4BrGSdj7wWJBKvq4ZG+/sPFlX+Y+pqRPZB2uRZYR
nGBwU7A6cmvxxmqNXL6cfq7pEtqiPakX8kxyXuKEH8PrIB2bKpiB/glQlozTVkLAhIX0qOhIA55B
ANYZ+3hh1JK6Cg07IDmXlYTIb0ffvzP/elckYxSbQeRXY3UU9AjThpxw0/PzxQa7A6K3gOoAvbKN
aQHqS1ybauqdvyPYQx0yz9Mdt4HPH3wNCNT7CJQ+1MZb0eELmJjnMjjRb0fZqT5YZbd8dyikgrb1
qF0cbooqAmY8r6+fjDwSgWWZdBzUn2OdlxSAQEjwWG6yeIx4zK5rPZZEVk47X6IE0O+IJ8EY9qt9
0w9bQ+dCO5evU5bD0K/hSXpXxVMtJxqv1vMX2vQaqe6rS0V7f7UtYyVNOqbIQ0hysRSE2vOjPS11
+7waO8JTFwmqHOHywX2UZpVYkWINv/xqAnWXqorwl9RB8f2NIIZ+LsQ7MjwZKbbtGdAH7BDm3drT
9aUj2VfqvLkHwwq3Jro6CaZ1b0hYrm8i9jKdujSpNN+3KOx1V0Q0LrSp2Fh4wb4Nxd/L8j8jETTF
zHScbGZS17zpYk8tshqsO5hU/lfWT1To2Jo2i1lWGdUa3+hujGaNcD5bwoxojhNx+NscgNFBOwgU
GYretmZooaHjpapacOO44QcACMTQ/3ovF8v5S2nAIwH17EaP5Go22RgyQld0qQxEFreayUbuaKO4
EIa+KK1XXgsNwr1C2vKHT8g3idxxAH6iNV79nbjH4L6l+xPb37jdHl0tqpcc5v9rJuZaCyDY+O2Q
xUSnYfbr7ywYDfVrG1/SUMims5z2XXPabNN1i2yeOK6UYi3gVdNU/xQ/HMlvJ59ATDFUDZD91Ku5
fmiuSfniHkgcaBBdmxffKt7T4fOIXEfAxSRGwHaNhfNwvlad95yrRjLK5viC/+adV7pz0dOGAsI/
Ft/z5kmjoUhChC4b/SQScjo5yG3hnbE+N3dGFDSY0RdhjSV5zNq/DvJV/7p9U1RlE9INVeVFPERJ
8k51vmYd58Ah3poUUYr0Q53sXh7PAyWEzYH0vx0cjoRp7A0RgIi56/JhGtgg0bJK8f2X4OHMhkjj
lURuNmKmgW4JcV9VOjDSCZjFUOisXzzsL1p18nfRwBbawy6OxWZM4i7GXK/p9OflHsXCCUimvYnK
zszkCzz3/Ynn/c7E8m7qeMRxIbEzaPF/dv+ic+0i7nuFWjWCRgZ28WBKa6PFvZoBDI3joZqw5s31
3kYCtWHCElWNm7Y71P8crgVPZ1xS5Qjbk/hewJGOO9kHiN9jszelNiIaNQqNevJmBDgfSsxyak9V
ofF5aIaLkKrXH7uzXUdb7H90AJy00Pu2FwHuk2z0RNISqTRqRWN7iCCooJNqq6hJkwDUSbOvuZRt
efBiPxkDu0UaSaDT0snDD9xu0dALqLDGQfY6GeLUYqulBffJyAcMXnXhKzRM3lWAkmZteAEoJA2+
z2UhMDjQ4Ve17rBWxyK4Vi6qjI0BgiStRNmm3G627UmOZ/5gwEj/fhdU9woE6tojbnrX7boSXPxx
AR5PnPZrFek1APcY5irU2HeSWkobKNlBEBqubTlOjZyAqEzUyhieOdC7ATV/fdaK+O5X8uE3L7aZ
Azdfnpu2KWrx090c9C2sKKmthzDT+Dayp/7UT6sAl7aHafGa60ty5j2cEgIs7GxiwP67KsDgbNlh
YyM5djVs+F77Hl0J5WPAUSiovKYPpM9JO+szapNxgGlF6r9Syrrjq0d9TSyb8YBSRu9mHMAw1ULg
T/Ex2mPKG356s2dVNV/04vI9ZBs2/4UJVmMdNmUwZTxxvoUIOsC3PNnCXu133Y1xhbhJh7zB++Jg
xkw+nwpmn5xSJ63rUv0g+xZXXUk/rJGGbj+FqqCsn7vh8gUiWZfd6p+TT/6Xa+mIjB88XdEx9hS4
eFk27EWCBfj5LxJgRuq8RCnQiD4JG89VIvhV1f9e4XTmL1s1A1H5Kq9HVASBx0XbK+7YVN105bgA
4V/xXKPa7UNl2Pdk2hgqDEKRAf3nsmRuIkD5/9elBLSV6AgIiivHsnmtKbNJlZn2Dj51p2Hk92Pa
tYggsF7uZsZe4+MpTechXcFF9bZhIqBNaWISkWQoU2EL9x3F2slGWentolZoRMjCGkQPGNeaINcB
DYReKxln72f9yXwHOUNu7ogq7C9knPsdB4XO8lX+YMcg+95IS4CX34f9uEjetDIFIV2ErQSOv0Tc
VZvnBGexJz8wlpafyCIYzctDyXmPZQs7MHTJPhk6gsOb3lVHAos8bRfj36WPWb11Z+JS/gEBfSmI
iNKfum8TTY6E21xX73v9ET9h4tKUcByGpwe04mzs0k5pbyPppCrBRWYVUwIe0u+De8AARme9o5cX
2zSPbMhqfqWP0G4DYEbSystCfQkLD1LCTvWFmJmItYMJtEFj62KnqmOCNHOesGqFR+J1Kttp2cBQ
4/+D8FNtT55aqVGsqwRaFhSnhiDFq1XAWQgdlZ1IRhGSa17X+Ao+VHO3UYXOgdbynZyjNLWfWZTZ
4+Fr8U6TGiGVUt2mUFQhvyUVs3cUoVxDe8skNBIerCUEmPNBiSK+rx2eeCFB3b1aiy6RJoDARILX
/4YZ3MNZWtvejA==
`protect end_protected
